module division (
	input logic [31:0] i_dividend, i_divisor,
	output logic [31:0] o_quotient,
	output logic [31:0] o_remainder
);



endmodule
