module reg0_32bit (
	output logic [31:0] RD
);

assign RD = 32'h0000_0000;

endmodule : reg0_32bit
	