/*
==================================================================================================
						  ____            _             _   _   _       _ _   
						 / ___|___  _ __ | |_ _ __ ___ | | | | | |_ __ (_) |_ 
						| |   / _ \| '_ \| __| '__/ _ \| | | | | | '_ \| | __|
						| |__| (_) | | | | |_| | | (_) | | | |_| | | | | | |_ 
						 \____\___/|_| |_|\__|_|  \___/|_|  \___/|_| |_|_|\__|
																						 
==================================================================================================
*/
module control_unit
(

);


endmodule 



/*
==================================================================================================
						  ___       _                          ____ _        _ 
						 |_ _|_ __ | |_ ___  __ _  ___ _ __   / ___| |_ _ __| |
						  | || '_ \| __/ _ \/ _` |/ _ \ '__| | |   | __| '__| |
						  | || | | | ||  __/ (_| |  __/ |    | |___| |_| |  | |
						 |___|_| |_|\__\___|\__, |\___|_|     \____|\__|_|  |_|
												  |___/                              
==================================================================================================
*/
module integer_ctrl
(

);


endmodule 


/*
==================================================================================================
	  __  __       _ _   _       _          ______  _       _     _         ____ _        _ 
	 |  \/  |_   _| | |_(_)_ __ | |_   _   / /  _ \(_)_   _(_) __| | ___   / ___| |_ _ __| |
	 | |\/| | | | | | __| | '_ \| | | | | / /| | | | \ \ / / |/ _` |/ _ \ | |   | __| '__| |
	 | |  | | |_| | | |_| | |_) | | |_| |/ / | |_| | |\ V /| | (_| |  __/ | |___| |_| |  | |
	 |_|  |_|\__,_|_|\__|_| .__/|_|\__, /_/  |____/|_| \_/ |_|\__,_|\___|  \____|\__|_|  |_|
								 |_|      |___/                                                    
==================================================================================================
*/
module mult_ctrl
(

);


endmodule 


/*
==================================================================================================
		  _____ _             _   _               ____       _       _      ____ _        _ 
		 |  ___| | ___   __ _| |_(_)_ __   __ _  |  _ \ ___ (_)_ __ | |_   / ___| |_ _ __| |
		 | |_  | |/ _ \ / _` | __| | '_ \ / _` | | |_) / _ \| | '_ \| __| | |   | __| '__| |
		 |  _| | | (_) | (_| | |_| | | | | (_| | |  __/ (_) | | | | | |_  | |___| |_| |  | |
		 |_|   |_|\___/ \__,_|\__|_|_| |_|\__, | |_|   \___/|_|_| |_|\__|  \____|\__|_|  |_|
													 |___/                                             
==================================================================================================
*/
module fp_ctrl
(

);


endmodule 


