module division (
	input logic [31:0] i_dividend, i_divisor,
	output logic [31:0] o_quotient,
	output logic [31:0] o_remainder
);

logic [30:0] result0, cout0;
logic [30:0] result1, cout1;
logic [30:0] result2, cout2;
logic [30:0] result3, cout3;
logic [30:0] result4, cout4;
logic [30:0] result5, cout5;
logic [30:0] result6, cout6;
logic [30:0] result7, cout7;
logic [30:0] result8, cout8;
logic [30:0] result9, cout9;
logic [30:0] result10, cout10;
logic [30:0] result11, cout11;
logic [30:0] result12, cout12;
logic [30:0] result13, cout13;
logic [30:0] result14, cout14;
logic [30:0] result15, cout15;
logic [30:0] result16, cout16;
logic [30:0] result17, cout17;
logic [30:0] result18, cout18;
logic [30:0] result19, cout19;
logic [30:0] result20, cout20;
logic [30:0] result21, cout21;
logic [30:0] result22, cout22;
logic [30:0] result23, cout23;
logic [30:0] result24, cout24;
logic [30:0] result25, cout25;
logic [30:0] result26, cout26;
logic [30:0] result27, cout27;
logic [30:0] result28, cout28;
logic [30:0] result29, cout29;
logic [30:0] result30, cout30;
logic [30:0] cout31;
logic [31:0] result31;
logic [31:0] quotient;

// Row 0
pu pu0_0 (.i_a(i_dividend[31]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[31]),
	 	   .o_result(result0[0]), .o_cout(cout0[0]));
pu pu0_1 (.i_a(0), .i_b(~i_divisor[1]), .i_cin(cout0[0]), .i_carry_output(quotient[31]),
	  	   .o_result(result0[1]), .o_cout(cout0[1]));
pu pu0_2 (.i_a(0), .i_b(~i_divisor[2]), .i_cin(cout0[1]), .i_carry_output(quotient[31]),
		   .o_result(result0[2]), .o_cout(cout0[2]));
pu pu0_3 (.i_a(0), .i_b(~i_divisor[3]), .i_cin(cout0[2]), .i_carry_output(quotient[31]),
		   .o_result(result0[3]), .o_cout(cout0[3]));
pu pu0_4 (.i_a(0), .i_b(~i_divisor[4]), .i_cin(cout0[3]), .i_carry_output(quotient[31]),
		   .o_result(result0[4]), .o_cout(cout0[4]));	
pu pu0_5 (.i_a(0), .i_b(~i_divisor[5]), .i_cin(cout0[4]), .i_carry_output(quotient[31]),
		   .o_result(result0[5]), .o_cout(cout0[5]));		  
pu pu0_6 (.i_a(0), .i_b(~i_divisor[6]), .i_cin(cout0[5]), .i_carry_output(quotient[31]),
		   .o_result(result0[6]), .o_cout(cout0[6]));			  
pu pu0_7 (.i_a(0), .i_b(~i_divisor[7]), .i_cin(cout0[6]), .i_carry_output(quotient[31]),
	 	   .o_result(result0[7]), .o_cout(cout0[7]));				  
pu pu0_8 (.i_a(0), .i_b(~i_divisor[8]), .i_cin(cout0[7]), .i_carry_output(quotient[31]),
         .o_result(result0[8]), .o_cout(cout0[8]));
pu pu0_9 (.i_a(0), .i_b(~i_divisor[9]), .i_cin(cout0[8]), .i_carry_output(quotient[31]),
         .o_result(result0[9]), .o_cout(cout0[9]));
pu pu0_10 (.i_a(0), .i_b(~i_divisor[10]), .i_cin(cout0[9]), .i_carry_output(quotient[31]),
          .o_result(result0[10]), .o_cout(cout0[10]));
pu pu0_11 (.i_a(0), .i_b(~i_divisor[11]), .i_cin(cout0[10]), .i_carry_output(quotient[31]),
          .o_result(result0[11]), .o_cout(cout0[11]));
pu pu0_12 (.i_a(0), .i_b(~i_divisor[12]), .i_cin(cout0[11]), .i_carry_output(quotient[31]),
          .o_result(result0[12]), .o_cout(cout0[12]));
pu pu0_13 (.i_a(0), .i_b(~i_divisor[13]), .i_cin(cout0[12]), .i_carry_output(quotient[31]),
          .o_result(result0[13]), .o_cout(cout0[13]));
pu pu0_14 (.i_a(0), .i_b(~i_divisor[14]), .i_cin(cout0[13]), .i_carry_output(quotient[31]),
          .o_result(result0[14]), .o_cout(cout0[14]));
pu pu0_15 (.i_a(0), .i_b(~i_divisor[15]), .i_cin(cout0[14]), .i_carry_output(quotient[31]),
          .o_result(result0[15]), .o_cout(cout0[15]));
pu pu0_16 (.i_a(0), .i_b(~i_divisor[16]), .i_cin(cout0[15]), .i_carry_output(quotient[31]),
          .o_result(result0[16]), .o_cout(cout0[16]));
pu pu0_17 (.i_a(0), .i_b(~i_divisor[17]), .i_cin(cout0[16]), .i_carry_output(quotient[31]),
          .o_result(result0[17]), .o_cout(cout0[17]));
pu pu0_18 (.i_a(0), .i_b(~i_divisor[18]), .i_cin(cout0[17]), .i_carry_output(quotient[31]),
          .o_result(result0[18]), .o_cout(cout0[18]));
pu pu0_19 (.i_a(0), .i_b(~i_divisor[19]), .i_cin(cout0[18]), .i_carry_output(quotient[31]),
          .o_result(result0[19]), .o_cout(cout0[19]));
pu pu0_20 (.i_a(0), .i_b(~i_divisor[20]), .i_cin(cout0[19]), .i_carry_output(quotient[31]),
          .o_result(result0[20]), .o_cout(cout0[20]));
pu pu0_21 (.i_a(0), .i_b(~i_divisor[21]), .i_cin(cout0[20]), .i_carry_output(quotient[31]),
          .o_result(result0[21]), .o_cout(cout0[21]));
pu pu0_22 (.i_a(0), .i_b(~i_divisor[22]), .i_cin(cout0[21]), .i_carry_output(quotient[31]),
          .o_result(result0[22]), .o_cout(cout0[22]));
pu pu0_23 (.i_a(0), .i_b(~i_divisor[23]), .i_cin(cout0[22]), .i_carry_output(quotient[31]),
          .o_result(result0[23]), .o_cout(cout0[23]));
pu pu0_24 (.i_a(0), .i_b(~i_divisor[24]), .i_cin(cout0[23]), .i_carry_output(quotient[31]),
          .o_result(result0[24]), .o_cout(cout0[24]));
pu pu0_25 (.i_a(0), .i_b(~i_divisor[25]), .i_cin(cout0[24]), .i_carry_output(quotient[31]),
          .o_result(result0[25]), .o_cout(cout0[25]));
pu pu0_26 (.i_a(0), .i_b(~i_divisor[26]), .i_cin(cout0[25]), .i_carry_output(quotient[31]),
          .o_result(result0[26]), .o_cout(cout0[26]));
pu pu0_27 (.i_a(0), .i_b(~i_divisor[27]), .i_cin(cout0[26]), .i_carry_output(quotient[31]),
          .o_result(result0[27]), .o_cout(cout0[27]));
pu pu0_28 (.i_a(0), .i_b(~i_divisor[28]), .i_cin(cout0[27]), .i_carry_output(quotient[31]),
          .o_result(result0[28]), .o_cout(cout0[28]));
pu pu0_29 (.i_a(0), .i_b(~i_divisor[29]), .i_cin(cout0[28]), .i_carry_output(quotient[31]),
          .o_result(result0[29]), .o_cout(cout0[29]));
pu pu0_30 (.i_a(0), .i_b(~i_divisor[30]), .i_cin(cout0[29]), .i_carry_output(quotient[31]),
          .o_result(result0[30]), .o_cout(cout0[30]));
pu pu0_31 (.i_a(0), .i_b(~i_divisor[31]), .i_cin(cout0[30]), .i_carry_output(quotient[31]),
          .o_cout(quotient[31]));

// Row 1
pu pu1_0 (.i_a(i_dividend[30]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[30]),
         .o_result(result1[0]), .o_cout(cout1[0]));
pu pu1_1 (.i_a(result0[0]), .i_b(~i_divisor[1]), .i_cin(cout1[0]), .i_carry_output(quotient[30]),
	  	   .o_result(result1[1]), .o_cout(cout1[1]));
pu pu1_2 (.i_a(result0[1]), .i_b(~i_divisor[2]), .i_cin(cout1[1]), .i_carry_output(quotient[30]),
	  	   .o_result(result1[2]), .o_cout(cout1[2]));
pu pu1_3 (.i_a(result0[2]), .i_b(~i_divisor[3]), .i_cin(cout1[2]), .i_carry_output(quotient[30]),
		   .o_result(result1[3]), .o_cout(cout1[3]));
pu pu1_4 (.i_a(result0[3]), .i_b(~i_divisor[4]), .i_cin(cout1[3]), .i_carry_output(quotient[30]),
		   .o_result(result1[4]), .o_cout(cout1[4]));
pu pu1_5 (.i_a(result0[4]), .i_b(~i_divisor[5]), .i_cin(cout1[4]), .i_carry_output(quotient[30]),
		   .o_result(result1[5]), .o_cout(cout1[5]));
pu pu1_6 (.i_a(result0[5]), .i_b(~i_divisor[6]), .i_cin(cout1[5]), .i_carry_output(quotient[30]),
		   .o_result(result1[6]), .o_cout(cout1[6]));
pu pu1_7 (.i_a(result0[6]), .i_b(~i_divisor[7]), .i_cin(cout1[6]), .i_carry_output(quotient[30]),
		   .o_result(result1[7]), .o_cout(cout1[7]));
pu pu1_8 (.i_a(result0[7]), .i_b(~i_divisor[8]), .i_cin(cout1[7]), .i_carry_output(quotient[30]),
		   .o_result(result1[8]), .o_cout(cout1[8]));
pu pu1_9 (.i_a(result0[8]), .i_b(~i_divisor[9]), .i_cin(cout1[8]), .i_carry_output(quotient[30]),
		   .o_result(result1[9]), .o_cout(cout1[9]));
pu pu1_10 (.i_a(result0[9]), .i_b(~i_divisor[10]), .i_cin(cout1[9]), .i_carry_output(quotient[30]),
		    .o_result(result1[10]), .o_cout(cout1[10]));
pu pu1_11 (.i_a(result0[10]), .i_b(~i_divisor[11]), .i_cin(cout1[10]), .i_carry_output(quotient[30]),
		    .o_result(result1[11]), .o_cout(cout1[11]));
pu pu1_12 (.i_a(result0[11]), .i_b(~i_divisor[12]), .i_cin(cout1[11]), .i_carry_output(quotient[30]),
		    .o_result(result1[12]), .o_cout(cout1[12]));
pu pu1_13 (.i_a(result0[12]), .i_b(~i_divisor[13]), .i_cin(cout1[12]), .i_carry_output(quotient[30]),
		    .o_result(result1[13]), .o_cout(cout1[13]));
pu pu1_14 (.i_a(result0[13]), .i_b(~i_divisor[14]), .i_cin(cout1[13]), .i_carry_output(quotient[30]),
		    .o_result(result1[14]), .o_cout(cout1[14]));
pu pu1_15 (.i_a(result0[14]), .i_b(~i_divisor[15]), .i_cin(cout1[14]), .i_carry_output(quotient[30]),
		    .o_result(result1[15]), .o_cout(cout1[15]));
pu pu1_16 (.i_a(result0[15]), .i_b(~i_divisor[16]), .i_cin(cout1[15]), .i_carry_output(quotient[30]),
		    .o_result(result1[16]), .o_cout(cout1[16]));
pu pu1_17 (.i_a(result0[16]), .i_b(~i_divisor[17]), .i_cin(cout1[16]), .i_carry_output(quotient[30]),
		    .o_result(result1[17]), .o_cout(cout1[17]));
pu pu1_18 (.i_a(result0[17]), .i_b(~i_divisor[18]), .i_cin(cout1[17]), .i_carry_output(quotient[30]),
		    .o_result(result1[18]), .o_cout(cout1[18]));
pu pu1_19 (.i_a(result0[18]), .i_b(~i_divisor[19]), .i_cin(cout1[18]), .i_carry_output(quotient[30]),
		    .o_result(result1[19]), .o_cout(cout1[19]));
pu pu1_20 (.i_a(result0[19]), .i_b(~i_divisor[20]), .i_cin(cout1[19]), .i_carry_output(quotient[30]),
		    .o_result(result1[20]), .o_cout(cout1[20]));
pu pu1_21 (.i_a(result0[20]), .i_b(~i_divisor[21]), .i_cin(cout1[20]), .i_carry_output(quotient[30]),
		    .o_result(result1[21]), .o_cout(cout1[21]));
pu pu1_22 (.i_a(result0[21]), .i_b(~i_divisor[22]), .i_cin(cout1[21]), .i_carry_output(quotient[30]),
		    .o_result(result1[22]), .o_cout(cout1[22]));
pu pu1_23 (.i_a(result0[22]), .i_b(~i_divisor[23]), .i_cin(cout1[22]), .i_carry_output(quotient[30]),
		    .o_result(result1[23]), .o_cout(cout1[23]));
pu pu1_24 (.i_a(result0[23]), .i_b(~i_divisor[24]), .i_cin(cout1[23]), .i_carry_output(quotient[30]),
		    .o_result(result1[24]), .o_cout(cout1[24]));
pu pu1_25 (.i_a(result0[24]), .i_b(~i_divisor[25]), .i_cin(cout1[24]), .i_carry_output(quotient[30]),
		    .o_result(result1[25]), .o_cout(cout1[25]));
pu pu1_26 (.i_a(result0[25]), .i_b(~i_divisor[26]), .i_cin(cout1[25]), .i_carry_output(quotient[30]),
		    .o_result(result1[26]), .o_cout(cout1[26]));
pu pu1_27 (.i_a(result0[26]), .i_b(~i_divisor[27]), .i_cin(cout1[26]), .i_carry_output(quotient[30]),
		    .o_result(result1[27]), .o_cout(cout1[27]));
pu pu1_28 (.i_a(result0[27]), .i_b(~i_divisor[28]), .i_cin(cout1[27]), .i_carry_output(quotient[30]),
		    .o_result(result1[28]), .o_cout(cout1[28]));
pu pu1_29 (.i_a(result0[28]), .i_b(~i_divisor[29]), .i_cin(cout1[28]), .i_carry_output(quotient[30]),
		    .o_result(result1[29]), .o_cout(cout1[29]));
pu pu1_30 (.i_a(result0[29]), .i_b(~i_divisor[30]), .i_cin(cout1[29]), .i_carry_output(quotient[30]),
		    .o_result(result1[30]), .o_cout(cout1[30]));
pu pu1_31 (.i_a(result0[30]), .i_b(~i_divisor[31]), .i_cin(cout1[30]), .i_carry_output(quotient[30]),
		    .o_cout(quotient[30]));

// Row 2
pu pu2_0 (.i_a(i_dividend[29]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[29]),
         .o_result(result2[0]), .o_cout(cout2[0]));			 
pu pu2_1 (.i_a(result1[0]), .i_b(~i_divisor[1]), .i_cin(cout2[0]), .i_carry_output(quotient[29]),
		.o_result(result2[1]), .o_cout(cout2[1]));
pu pu2_2 (.i_a(result1[1]), .i_b(~i_divisor[2]), .i_cin(cout2[1]), .i_carry_output(quotient[29]),
		.o_result(result2[2]), .o_cout(cout2[2]));
pu pu2_3 (.i_a(result1[2]), .i_b(~i_divisor[3]), .i_cin(cout2[2]), .i_carry_output(quotient[29]),
		.o_result(result2[3]), .o_cout(cout2[3]));
pu pu2_4 (.i_a(result1[3]), .i_b(~i_divisor[4]), .i_cin(cout2[3]), .i_carry_output(quotient[29]),
		.o_result(result2[4]), .o_cout(cout2[4]));
pu pu2_5 (.i_a(result1[4]), .i_b(~i_divisor[5]), .i_cin(cout2[4]), .i_carry_output(quotient[29]),
		.o_result(result2[5]), .o_cout(cout2[5]));
pu pu2_6 (.i_a(result1[5]), .i_b(~i_divisor[6]), .i_cin(cout2[5]), .i_carry_output(quotient[29]),
		.o_result(result2[6]), .o_cout(cout2[6]));
pu pu2_7 (.i_a(result1[6]), .i_b(~i_divisor[7]), .i_cin(cout2[6]), .i_carry_output(quotient[29]),
		.o_result(result2[7]), .o_cout(cout2[7]));
pu pu2_8 (.i_a(result1[7]), .i_b(~i_divisor[8]), .i_cin(cout2[7]), .i_carry_output(quotient[29]),
		.o_result(result2[8]), .o_cout(cout2[8]));
pu pu2_9 (.i_a(result1[8]), .i_b(~i_divisor[9]), .i_cin(cout2[8]), .i_carry_output(quotient[29]),
		.o_result(result2[9]), .o_cout(cout2[9]));
pu pu2_10 (.i_a(result1[9]), .i_b(~i_divisor[10]), .i_cin(cout2[9]), .i_carry_output(quotient[29]),
		.o_result(result2[10]), .o_cout(cout2[10]));
pu pu2_11 (.i_a(result1[10]), .i_b(~i_divisor[11]), .i_cin(cout2[10]), .i_carry_output(quotient[29]),
		.o_result(result2[11]), .o_cout(cout2[11]));
pu pu2_12 (.i_a(result1[11]), .i_b(~i_divisor[12]), .i_cin(cout2[11]), .i_carry_output(quotient[29]),
		.o_result(result2[12]), .o_cout(cout2[12]));
pu pu2_13 (.i_a(result1[12]), .i_b(~i_divisor[13]), .i_cin(cout2[12]), .i_carry_output(quotient[29]),
		.o_result(result2[13]), .o_cout(cout2[13]));
pu pu2_14 (.i_a(result1[13]), .i_b(~i_divisor[14]), .i_cin(cout2[13]), .i_carry_output(quotient[29]),
		.o_result(result2[14]), .o_cout(cout2[14]));
pu pu2_15 (.i_a(result1[14]), .i_b(~i_divisor[15]), .i_cin(cout2[14]), .i_carry_output(quotient[29]),
		.o_result(result2[15]), .o_cout(cout2[15]));
pu pu2_16 (.i_a(result1[15]), .i_b(~i_divisor[16]), .i_cin(cout2[15]), .i_carry_output(quotient[29]),
		.o_result(result2[16]), .o_cout(cout2[16]));
pu pu2_17 (.i_a(result1[16]), .i_b(~i_divisor[17]), .i_cin(cout2[16]), .i_carry_output(quotient[29]),
		.o_result(result2[17]), .o_cout(cout2[17]));
pu pu2_18 (.i_a(result1[17]), .i_b(~i_divisor[18]), .i_cin(cout2[17]), .i_carry_output(quotient[29]),
		.o_result(result2[18]), .o_cout(cout2[18]));
pu pu2_19 (.i_a(result1[18]), .i_b(~i_divisor[19]), .i_cin(cout2[18]), .i_carry_output(quotient[29]),
		.o_result(result2[19]), .o_cout(cout2[19]));
pu pu2_20 (.i_a(result1[19]), .i_b(~i_divisor[20]), .i_cin(cout2[19]), .i_carry_output(quotient[29]),
		.o_result(result2[20]), .o_cout(cout2[20]));
pu pu2_21 (.i_a(result1[20]), .i_b(~i_divisor[21]), .i_cin(cout2[20]), .i_carry_output(quotient[29]),
		.o_result(result2[21]), .o_cout(cout2[21]));
pu pu2_22 (.i_a(result1[21]), .i_b(~i_divisor[22]), .i_cin(cout2[21]), .i_carry_output(quotient[29]),
		.o_result(result2[22]), .o_cout(cout2[22]));
pu pu2_23 (.i_a(result1[22]), .i_b(~i_divisor[23]), .i_cin(cout2[22]), .i_carry_output(quotient[29]),
		.o_result(result2[23]), .o_cout(cout2[23]));
pu pu2_24 (.i_a(result1[23]), .i_b(~i_divisor[24]), .i_cin(cout2[23]), .i_carry_output(quotient[29]),
		.o_result(result2[24]), .o_cout(cout2[24]));
pu pu2_25 (.i_a(result1[24]), .i_b(~i_divisor[25]), .i_cin(cout2[24]), .i_carry_output(quotient[29]),
		.o_result(result2[25]), .o_cout(cout2[25]));
pu pu2_26 (.i_a(result1[25]), .i_b(~i_divisor[26]), .i_cin(cout2[25]), .i_carry_output(quotient[29]),
		.o_result(result2[26]), .o_cout(cout2[26]));
pu pu2_27 (.i_a(result1[26]), .i_b(~i_divisor[27]), .i_cin(cout2[26]), .i_carry_output(quotient[29]),
		.o_result(result2[27]), .o_cout(cout2[27]));
pu pu2_28 (.i_a(result1[27]), .i_b(~i_divisor[28]), .i_cin(cout2[27]), .i_carry_output(quotient[29]),
		.o_result(result2[28]), .o_cout(cout2[28]));
pu pu2_29 (.i_a(result1[28]), .i_b(~i_divisor[29]), .i_cin(cout2[28]), .i_carry_output(quotient[29]),
		.o_result(result2[29]), .o_cout(cout2[29]));
pu pu2_30 (.i_a(result1[29]), .i_b(~i_divisor[30]), .i_cin(cout2[29]), .i_carry_output(quotient[29]),
		.o_result(result2[30]), .o_cout(cout2[30]));
pu pu2_31 (.i_a(result1[30]), .i_b(~i_divisor[31]), .i_cin(cout2[30]), .i_carry_output(quotient[29]),
		.o_cout(quotient[29]));

// Row 3	
pu pu3_0 (.i_a(i_dividend[28]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[28]),
         .o_result(result3[0]), .o_cout(cout3[0]));		
pu pu3_1 (.i_a(result2[0]), .i_b(~i_divisor[1]), .i_cin(cout3[0]), .i_carry_output(quotient[28]),
		.o_result(result3[1]), .o_cout(cout3[1]));
pu pu3_2 (.i_a(result2[1]), .i_b(~i_divisor[2]), .i_cin(cout3[1]), .i_carry_output(quotient[28]),
		.o_result(result3[2]), .o_cout(cout3[2]));
pu pu3_3 (.i_a(result2[2]), .i_b(~i_divisor[3]), .i_cin(cout3[2]), .i_carry_output(quotient[28]),
		.o_result(result3[3]), .o_cout(cout3[3]));
pu pu3_4 (.i_a(result2[3]), .i_b(~i_divisor[4]), .i_cin(cout3[3]), .i_carry_output(quotient[28]),
		.o_result(result3[4]), .o_cout(cout3[4]));
pu pu3_5 (.i_a(result2[4]), .i_b(~i_divisor[5]), .i_cin(cout3[4]), .i_carry_output(quotient[28]),
		.o_result(result3[5]), .o_cout(cout3[5]));
pu pu3_6 (.i_a(result2[5]), .i_b(~i_divisor[6]), .i_cin(cout3[5]), .i_carry_output(quotient[28]),
		.o_result(result3[6]), .o_cout(cout3[6]));
pu pu3_7 (.i_a(result2[6]), .i_b(~i_divisor[7]), .i_cin(cout3[6]), .i_carry_output(quotient[28]),
		.o_result(result3[7]), .o_cout(cout3[7]));
pu pu3_8 (.i_a(result2[7]), .i_b(~i_divisor[8]), .i_cin(cout3[7]), .i_carry_output(quotient[28]),
		.o_result(result3[8]), .o_cout(cout3[8]));
pu pu3_9 (.i_a(result2[8]), .i_b(~i_divisor[9]), .i_cin(cout3[8]), .i_carry_output(quotient[28]),
		.o_result(result3[9]), .o_cout(cout3[9]));
pu pu3_10 (.i_a(result2[9]), .i_b(~i_divisor[10]), .i_cin(cout3[9]), .i_carry_output(quotient[28]),
		.o_result(result3[10]), .o_cout(cout3[10]));
pu pu3_11 (.i_a(result2[10]), .i_b(~i_divisor[11]), .i_cin(cout3[10]), .i_carry_output(quotient[28]),
		.o_result(result3[11]), .o_cout(cout3[11]));
pu pu3_12 (.i_a(result2[11]), .i_b(~i_divisor[12]), .i_cin(cout3[11]), .i_carry_output(quotient[28]),
		.o_result(result3[12]), .o_cout(cout3[12]));
pu pu3_13 (.i_a(result2[12]), .i_b(~i_divisor[13]), .i_cin(cout3[12]), .i_carry_output(quotient[28]),
		.o_result(result3[13]), .o_cout(cout3[13]));
pu pu3_14 (.i_a(result2[13]), .i_b(~i_divisor[14]), .i_cin(cout3[13]), .i_carry_output(quotient[28]),
		.o_result(result3[14]), .o_cout(cout3[14]));
pu pu3_15 (.i_a(result2[14]), .i_b(~i_divisor[15]), .i_cin(cout3[14]), .i_carry_output(quotient[28]),
		.o_result(result3[15]), .o_cout(cout3[15]));
pu pu3_16 (.i_a(result2[15]), .i_b(~i_divisor[16]), .i_cin(cout3[15]), .i_carry_output(quotient[28]),
		.o_result(result3[16]), .o_cout(cout3[16]));
pu pu3_17 (.i_a(result2[16]), .i_b(~i_divisor[17]), .i_cin(cout3[16]), .i_carry_output(quotient[28]),
		.o_result(result3[17]), .o_cout(cout3[17]));
pu pu3_18 (.i_a(result2[17]), .i_b(~i_divisor[18]), .i_cin(cout3[17]), .i_carry_output(quotient[28]),
		.o_result(result3[18]), .o_cout(cout3[18]));
pu pu3_19 (.i_a(result2[18]), .i_b(~i_divisor[19]), .i_cin(cout3[18]), .i_carry_output(quotient[28]),
		.o_result(result3[19]), .o_cout(cout3[19]));
pu pu3_20 (.i_a(result2[19]), .i_b(~i_divisor[20]), .i_cin(cout3[19]), .i_carry_output(quotient[28]),
		.o_result(result3[20]), .o_cout(cout3[20]));
pu pu3_21 (.i_a(result2[20]), .i_b(~i_divisor[21]), .i_cin(cout3[20]), .i_carry_output(quotient[28]),
		.o_result(result3[21]), .o_cout(cout3[21]));
pu pu3_22 (.i_a(result2[21]), .i_b(~i_divisor[22]), .i_cin(cout3[21]), .i_carry_output(quotient[28]),
		.o_result(result3[22]), .o_cout(cout3[22]));
pu pu3_23 (.i_a(result2[22]), .i_b(~i_divisor[23]), .i_cin(cout3[22]), .i_carry_output(quotient[28]),
		.o_result(result3[23]), .o_cout(cout3[23]));
pu pu3_24 (.i_a(result2[23]), .i_b(~i_divisor[24]), .i_cin(cout3[23]), .i_carry_output(quotient[28]),
		.o_result(result3[24]), .o_cout(cout3[24]));
pu pu3_25 (.i_a(result2[24]), .i_b(~i_divisor[25]), .i_cin(cout3[24]), .i_carry_output(quotient[28]),
		.o_result(result3[25]), .o_cout(cout3[25]));
pu pu3_26 (.i_a(result2[25]), .i_b(~i_divisor[26]), .i_cin(cout3[25]), .i_carry_output(quotient[28]),
		.o_result(result3[26]), .o_cout(cout3[26]));
pu pu3_27 (.i_a(result2[26]), .i_b(~i_divisor[27]), .i_cin(cout3[26]), .i_carry_output(quotient[28]),
		.o_result(result3[27]), .o_cout(cout3[27]));
pu pu3_28 (.i_a(result2[27]), .i_b(~i_divisor[28]), .i_cin(cout3[27]), .i_carry_output(quotient[28]),
		.o_result(result3[28]), .o_cout(cout3[28]));
pu pu3_29 (.i_a(result2[28]), .i_b(~i_divisor[29]), .i_cin(cout3[28]), .i_carry_output(quotient[28]),
		.o_result(result3[29]), .o_cout(cout3[29]));
pu pu3_30 (.i_a(result2[29]), .i_b(~i_divisor[30]), .i_cin(cout3[29]), .i_carry_output(quotient[28]),
		.o_result(result3[30]), .o_cout(cout3[30]));
pu pu3_31 (.i_a(result2[30]), .i_b(~i_divisor[31]), .i_cin(cout3[30]), .i_carry_output(quotient[28]),
		.o_cout(quotient[28]));

// Row 4
pu pu4_0 (.i_a(i_dividend[27]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[27]),
         .o_result(result4[0]), .o_cout(cout4[0]));
pu pu4_1 (.i_a(result3[0]), .i_b(~i_divisor[1]), .i_cin(cout4[0]), .i_carry_output(quotient[27]),
		.o_result(result4[1]), .o_cout(cout4[1]));
pu pu4_2 (.i_a(result3[1]), .i_b(~i_divisor[2]), .i_cin(cout4[1]), .i_carry_output(quotient[27]),
		.o_result(result4[2]), .o_cout(cout4[2]));
pu pu4_3 (.i_a(result3[2]), .i_b(~i_divisor[3]), .i_cin(cout4[2]), .i_carry_output(quotient[27]),
		.o_result(result4[3]), .o_cout(cout4[3]));
pu pu4_4 (.i_a(result3[3]), .i_b(~i_divisor[4]), .i_cin(cout4[3]), .i_carry_output(quotient[27]),
		.o_result(result4[4]), .o_cout(cout4[4]));
pu pu4_5 (.i_a(result3[4]), .i_b(~i_divisor[5]), .i_cin(cout4[4]), .i_carry_output(quotient[27]),
		.o_result(result4[5]), .o_cout(cout4[5]));
pu pu4_6 (.i_a(result3[5]), .i_b(~i_divisor[6]), .i_cin(cout4[5]), .i_carry_output(quotient[27]),
		.o_result(result4[6]), .o_cout(cout4[6]));
pu pu4_7 (.i_a(result3[6]), .i_b(~i_divisor[7]), .i_cin(cout4[6]), .i_carry_output(quotient[27]),
		.o_result(result4[7]), .o_cout(cout4[7]));
pu pu4_8 (.i_a(result3[7]), .i_b(~i_divisor[8]), .i_cin(cout4[7]), .i_carry_output(quotient[27]),
		.o_result(result4[8]), .o_cout(cout4[8]));
pu pu4_9 (.i_a(result3[8]), .i_b(~i_divisor[9]), .i_cin(cout4[8]), .i_carry_output(quotient[27]),
		.o_result(result4[9]), .o_cout(cout4[9]));
pu pu4_10 (.i_a(result3[9]), .i_b(~i_divisor[10]), .i_cin(cout4[9]), .i_carry_output(quotient[27]),
		.o_result(result4[10]), .o_cout(cout4[10]));
pu pu4_11 (.i_a(result3[10]), .i_b(~i_divisor[11]), .i_cin(cout4[10]), .i_carry_output(quotient[27]),
		.o_result(result4[11]), .o_cout(cout4[11]));
pu pu4_12 (.i_a(result3[11]), .i_b(~i_divisor[12]), .i_cin(cout4[11]), .i_carry_output(quotient[27]),
		.o_result(result4[12]), .o_cout(cout4[12]));
pu pu4_13 (.i_a(result3[12]), .i_b(~i_divisor[13]), .i_cin(cout4[12]), .i_carry_output(quotient[27]),
		.o_result(result4[13]), .o_cout(cout4[13]));
pu pu4_14 (.i_a(result3[13]), .i_b(~i_divisor[14]), .i_cin(cout4[13]), .i_carry_output(quotient[27]),
		.o_result(result4[14]), .o_cout(cout4[14]));
pu pu4_15 (.i_a(result3[14]), .i_b(~i_divisor[15]), .i_cin(cout4[14]), .i_carry_output(quotient[27]),
		.o_result(result4[15]), .o_cout(cout4[15]));
pu pu4_16 (.i_a(result3[15]), .i_b(~i_divisor[16]), .i_cin(cout4[15]), .i_carry_output(quotient[27]),
		.o_result(result4[16]), .o_cout(cout4[16]));
pu pu4_17 (.i_a(result3[16]), .i_b(~i_divisor[17]), .i_cin(cout4[16]), .i_carry_output(quotient[27]),
		.o_result(result4[17]), .o_cout(cout4[17]));
pu pu4_18 (.i_a(result3[17]), .i_b(~i_divisor[18]), .i_cin(cout4[17]), .i_carry_output(quotient[27]),
		.o_result(result4[18]), .o_cout(cout4[18]));
pu pu4_19 (.i_a(result3[18]), .i_b(~i_divisor[19]), .i_cin(cout4[18]), .i_carry_output(quotient[27]),
		.o_result(result4[19]), .o_cout(cout4[19]));
pu pu4_20 (.i_a(result3[19]), .i_b(~i_divisor[20]), .i_cin(cout4[19]), .i_carry_output(quotient[27]),
		.o_result(result4[20]), .o_cout(cout4[20]));
pu pu4_21 (.i_a(result3[20]), .i_b(~i_divisor[21]), .i_cin(cout4[20]), .i_carry_output(quotient[27]),
		.o_result(result4[21]), .o_cout(cout4[21]));
pu pu4_22 (.i_a(result3[21]), .i_b(~i_divisor[22]), .i_cin(cout4[21]), .i_carry_output(quotient[27]),
		.o_result(result4[22]), .o_cout(cout4[22]));
pu pu4_23 (.i_a(result3[22]), .i_b(~i_divisor[23]), .i_cin(cout4[22]), .i_carry_output(quotient[27]),
		.o_result(result4[23]), .o_cout(cout4[23]));
pu pu4_24 (.i_a(result3[23]), .i_b(~i_divisor[24]), .i_cin(cout4[23]), .i_carry_output(quotient[27]),
		.o_result(result4[24]), .o_cout(cout4[24]));
pu pu4_25 (.i_a(result3[24]), .i_b(~i_divisor[25]), .i_cin(cout4[24]), .i_carry_output(quotient[27]),
		.o_result(result4[25]), .o_cout(cout4[25]));
pu pu4_26 (.i_a(result3[25]), .i_b(~i_divisor[26]), .i_cin(cout4[25]), .i_carry_output(quotient[27]),
		.o_result(result4[26]), .o_cout(cout4[26]));
pu pu4_27 (.i_a(result3[26]), .i_b(~i_divisor[27]), .i_cin(cout4[26]), .i_carry_output(quotient[27]),
		.o_result(result4[27]), .o_cout(cout4[27]));
pu pu4_28 (.i_a(result3[27]), .i_b(~i_divisor[28]), .i_cin(cout4[27]), .i_carry_output(quotient[27]),
		.o_result(result4[28]), .o_cout(cout4[28]));
pu pu4_29 (.i_a(result3[28]), .i_b(~i_divisor[29]), .i_cin(cout4[28]), .i_carry_output(quotient[27]),
		.o_result(result4[29]), .o_cout(cout4[29]));
pu pu4_30 (.i_a(result3[29]), .i_b(~i_divisor[30]), .i_cin(cout4[29]), .i_carry_output(quotient[27]),
		.o_result(result4[30]), .o_cout(cout4[30]));
pu pu4_31 (.i_a(result3[30]), .i_b(~i_divisor[31]), .i_cin(cout4[30]), .i_carry_output(quotient[27]),
		.o_cout(quotient[27]));

// Row 5
pu pu5_0 (.i_a(i_dividend[26]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[26]),
         .o_result(result5[0]), .o_cout(cout5[0]));
pu pu5_1 (.i_a(result4[0]), .i_b(~i_divisor[1]), .i_cin(cout5[0]), .i_carry_output(quotient[26]),
		.o_result(result5[1]), .o_cout(cout5[1]));
pu pu5_2 (.i_a(result4[1]), .i_b(~i_divisor[2]), .i_cin(cout5[1]), .i_carry_output(quotient[26]),
		.o_result(result5[2]), .o_cout(cout5[2]));
pu pu5_3 (.i_a(result4[2]), .i_b(~i_divisor[3]), .i_cin(cout5[2]), .i_carry_output(quotient[26]),
		.o_result(result5[3]), .o_cout(cout5[3]));
pu pu5_4 (.i_a(result4[3]), .i_b(~i_divisor[4]), .i_cin(cout5[3]), .i_carry_output(quotient[26]),
		.o_result(result5[4]), .o_cout(cout5[4]));
pu pu5_5 (.i_a(result4[4]), .i_b(~i_divisor[5]), .i_cin(cout5[4]), .i_carry_output(quotient[26]),
		.o_result(result5[5]), .o_cout(cout5[5]));
pu pu5_6 (.i_a(result4[5]), .i_b(~i_divisor[6]), .i_cin(cout5[5]), .i_carry_output(quotient[26]),
		.o_result(result5[6]), .o_cout(cout5[6]));
pu pu5_7 (.i_a(result4[6]), .i_b(~i_divisor[7]), .i_cin(cout5[6]), .i_carry_output(quotient[26]),
		.o_result(result5[7]), .o_cout(cout5[7]));
pu pu5_8 (.i_a(result4[7]), .i_b(~i_divisor[8]), .i_cin(cout5[7]), .i_carry_output(quotient[26]),
		.o_result(result5[8]), .o_cout(cout5[8]));
pu pu5_9 (.i_a(result4[8]), .i_b(~i_divisor[9]), .i_cin(cout5[8]), .i_carry_output(quotient[26]),
		.o_result(result5[9]), .o_cout(cout5[9]));
pu pu5_10 (.i_a(result4[9]), .i_b(~i_divisor[10]), .i_cin(cout5[9]), .i_carry_output(quotient[26]),
		.o_result(result5[10]), .o_cout(cout5[10]));
pu pu5_11 (.i_a(result4[10]), .i_b(~i_divisor[11]), .i_cin(cout5[10]), .i_carry_output(quotient[26]),
		.o_result(result5[11]), .o_cout(cout5[11]));
pu pu5_12 (.i_a(result4[11]), .i_b(~i_divisor[12]), .i_cin(cout5[11]), .i_carry_output(quotient[26]),
		.o_result(result5[12]), .o_cout(cout5[12]));
pu pu5_13 (.i_a(result4[12]), .i_b(~i_divisor[13]), .i_cin(cout5[12]), .i_carry_output(quotient[26]),
		.o_result(result5[13]), .o_cout(cout5[13]));
pu pu5_14 (.i_a(result4[13]), .i_b(~i_divisor[14]), .i_cin(cout5[13]), .i_carry_output(quotient[26]),
		.o_result(result5[14]), .o_cout(cout5[14]));
pu pu5_15 (.i_a(result4[14]), .i_b(~i_divisor[15]), .i_cin(cout5[14]), .i_carry_output(quotient[26]),
		.o_result(result5[15]), .o_cout(cout5[15]));
pu pu5_16 (.i_a(result4[15]), .i_b(~i_divisor[16]), .i_cin(cout5[15]), .i_carry_output(quotient[26]),
		.o_result(result5[16]), .o_cout(cout5[16]));
pu pu5_17 (.i_a(result4[16]), .i_b(~i_divisor[17]), .i_cin(cout5[16]), .i_carry_output(quotient[26]),
		.o_result(result5[17]), .o_cout(cout5[17]));
pu pu5_18 (.i_a(result4[17]), .i_b(~i_divisor[18]), .i_cin(cout5[17]), .i_carry_output(quotient[26]),
		.o_result(result5[18]), .o_cout(cout5[18]));
pu pu5_19 (.i_a(result4[18]), .i_b(~i_divisor[19]), .i_cin(cout5[18]), .i_carry_output(quotient[26]),
		.o_result(result5[19]), .o_cout(cout5[19]));
pu pu5_20 (.i_a(result4[19]), .i_b(~i_divisor[20]), .i_cin(cout5[19]), .i_carry_output(quotient[26]),
		.o_result(result5[20]), .o_cout(cout5[20]));
pu pu5_21 (.i_a(result4[20]), .i_b(~i_divisor[21]), .i_cin(cout5[20]), .i_carry_output(quotient[26]),
		.o_result(result5[21]), .o_cout(cout5[21]));
pu pu5_22 (.i_a(result4[21]), .i_b(~i_divisor[22]), .i_cin(cout5[21]), .i_carry_output(quotient[26]),
		.o_result(result5[22]), .o_cout(cout5[22]));
pu pu5_23 (.i_a(result4[22]), .i_b(~i_divisor[23]), .i_cin(cout5[22]), .i_carry_output(quotient[26]),
		.o_result(result5[23]), .o_cout(cout5[23]));
pu pu5_24 (.i_a(result4[23]), .i_b(~i_divisor[24]), .i_cin(cout5[23]), .i_carry_output(quotient[26]),
		.o_result(result5[24]), .o_cout(cout5[24]));
pu pu5_25 (.i_a(result4[24]), .i_b(~i_divisor[25]), .i_cin(cout5[24]), .i_carry_output(quotient[26]),
		.o_result(result5[25]), .o_cout(cout5[25]));
pu pu5_26 (.i_a(result4[25]), .i_b(~i_divisor[26]), .i_cin(cout5[25]), .i_carry_output(quotient[26]),
		.o_result(result5[26]), .o_cout(cout5[26]));
pu pu5_27 (.i_a(result4[26]), .i_b(~i_divisor[27]), .i_cin(cout5[26]), .i_carry_output(quotient[26]),
		.o_result(result5[27]), .o_cout(cout5[27]));
pu pu5_28 (.i_a(result4[27]), .i_b(~i_divisor[28]), .i_cin(cout5[27]), .i_carry_output(quotient[26]),
		.o_result(result5[28]), .o_cout(cout5[28]));
pu pu5_29 (.i_a(result4[28]), .i_b(~i_divisor[29]), .i_cin(cout5[28]), .i_carry_output(quotient[26]),
		.o_result(result5[29]), .o_cout(cout5[29]));
pu pu5_30 (.i_a(result4[29]), .i_b(~i_divisor[30]), .i_cin(cout5[29]), .i_carry_output(quotient[26]),
		.o_result(result5[30]), .o_cout(cout5[30]));
pu pu5_31 (.i_a(result4[30]), .i_b(~i_divisor[31]), .i_cin(cout5[30]), .i_carry_output(quotient[26]),
		.o_cout(quotient[26]));
	
// Row 6
pu pu6_0 (.i_a(i_dividend[25]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[25]),
         .o_result(result6[0]), .o_cout(cout6[0]));
pu pu6_1 (.i_a(result5[0]), .i_b(~i_divisor[1]), .i_cin(cout6[0]), .i_carry_output(quotient[25]),
		.o_result(result6[1]), .o_cout(cout6[1]));
pu pu6_2 (.i_a(result5[1]), .i_b(~i_divisor[2]), .i_cin(cout6[1]), .i_carry_output(quotient[25]),
		.o_result(result6[2]), .o_cout(cout6[2]));
pu pu6_3 (.i_a(result5[2]), .i_b(~i_divisor[3]), .i_cin(cout6[2]), .i_carry_output(quotient[25]),
		.o_result(result6[3]), .o_cout(cout6[3]));
pu pu6_4 (.i_a(result5[3]), .i_b(~i_divisor[4]), .i_cin(cout6[3]), .i_carry_output(quotient[25]),
		.o_result(result6[4]), .o_cout(cout6[4]));
pu pu6_5 (.i_a(result5[4]), .i_b(~i_divisor[5]), .i_cin(cout6[4]), .i_carry_output(quotient[25]),
		.o_result(result6[5]), .o_cout(cout6[5]));
pu pu6_6 (.i_a(result5[5]), .i_b(~i_divisor[6]), .i_cin(cout6[5]), .i_carry_output(quotient[25]),
		.o_result(result6[6]), .o_cout(cout6[6]));
pu pu6_7 (.i_a(result5[6]), .i_b(~i_divisor[7]), .i_cin(cout6[6]), .i_carry_output(quotient[25]),
		.o_result(result6[7]), .o_cout(cout6[7]));
pu pu6_8 (.i_a(result5[7]), .i_b(~i_divisor[8]), .i_cin(cout6[7]), .i_carry_output(quotient[25]),
		.o_result(result6[8]), .o_cout(cout6[8]));
pu pu6_9 (.i_a(result5[8]), .i_b(~i_divisor[9]), .i_cin(cout6[8]), .i_carry_output(quotient[25]),
		.o_result(result6[9]), .o_cout(cout6[9]));
pu pu6_10 (.i_a(result5[9]), .i_b(~i_divisor[10]), .i_cin(cout6[9]), .i_carry_output(quotient[25]),
		.o_result(result6[10]), .o_cout(cout6[10]));
pu pu6_11 (.i_a(result5[10]), .i_b(~i_divisor[11]), .i_cin(cout6[10]), .i_carry_output(quotient[25]),
		.o_result(result6[11]), .o_cout(cout6[11]));
pu pu6_12 (.i_a(result5[11]), .i_b(~i_divisor[12]), .i_cin(cout6[11]), .i_carry_output(quotient[25]),
		.o_result(result6[12]), .o_cout(cout6[12]));
pu pu6_13 (.i_a(result5[12]), .i_b(~i_divisor[13]), .i_cin(cout6[12]), .i_carry_output(quotient[25]),
		.o_result(result6[13]), .o_cout(cout6[13]));
pu pu6_14 (.i_a(result5[13]), .i_b(~i_divisor[14]), .i_cin(cout6[13]), .i_carry_output(quotient[25]),
		.o_result(result6[14]), .o_cout(cout6[14]));
pu pu6_15 (.i_a(result5[14]), .i_b(~i_divisor[15]), .i_cin(cout6[14]), .i_carry_output(quotient[25]),
		.o_result(result6[15]), .o_cout(cout6[15]));
pu pu6_16 (.i_a(result5[15]), .i_b(~i_divisor[16]), .i_cin(cout6[15]), .i_carry_output(quotient[25]),
		.o_result(result6[16]), .o_cout(cout6[16]));
pu pu6_17 (.i_a(result5[16]), .i_b(~i_divisor[17]), .i_cin(cout6[16]), .i_carry_output(quotient[25]),
		.o_result(result6[17]), .o_cout(cout6[17]));
pu pu6_18 (.i_a(result5[17]), .i_b(~i_divisor[18]), .i_cin(cout6[17]), .i_carry_output(quotient[25]),
		.o_result(result6[18]), .o_cout(cout6[18]));
pu pu6_19 (.i_a(result5[18]), .i_b(~i_divisor[19]), .i_cin(cout6[18]), .i_carry_output(quotient[25]),
		.o_result(result6[19]), .o_cout(cout6[19]));
pu pu6_20 (.i_a(result5[19]), .i_b(~i_divisor[20]), .i_cin(cout6[19]), .i_carry_output(quotient[25]),
		.o_result(result6[20]), .o_cout(cout6[20]));
pu pu6_21 (.i_a(result5[20]), .i_b(~i_divisor[21]), .i_cin(cout6[20]), .i_carry_output(quotient[25]),
		.o_result(result6[21]), .o_cout(cout6[21]));
pu pu6_22 (.i_a(result5[21]), .i_b(~i_divisor[22]), .i_cin(cout6[21]), .i_carry_output(quotient[25]),
		.o_result(result6[22]), .o_cout(cout6[22]));
pu pu6_23 (.i_a(result5[22]), .i_b(~i_divisor[23]), .i_cin(cout6[22]), .i_carry_output(quotient[25]),
		.o_result(result6[23]), .o_cout(cout6[23]));
pu pu6_24 (.i_a(result5[23]), .i_b(~i_divisor[24]), .i_cin(cout6[23]), .i_carry_output(quotient[25]),
		.o_result(result6[24]), .o_cout(cout6[24]));
pu pu6_25 (.i_a(result5[24]), .i_b(~i_divisor[25]), .i_cin(cout6[24]), .i_carry_output(quotient[25]),
		.o_result(result6[25]), .o_cout(cout6[25]));
pu pu6_26 (.i_a(result5[25]), .i_b(~i_divisor[26]), .i_cin(cout6[25]), .i_carry_output(quotient[25]),
		.o_result(result6[26]), .o_cout(cout6[26]));
pu pu6_27 (.i_a(result5[26]), .i_b(~i_divisor[27]), .i_cin(cout6[26]), .i_carry_output(quotient[25]),
		.o_result(result6[27]), .o_cout(cout6[27]));
pu pu6_28 (.i_a(result5[27]), .i_b(~i_divisor[28]), .i_cin(cout6[27]), .i_carry_output(quotient[25]),
		.o_result(result6[28]), .o_cout(cout6[28]));
pu pu6_29 (.i_a(result5[28]), .i_b(~i_divisor[29]), .i_cin(cout6[28]), .i_carry_output(quotient[25]),
		.o_result(result6[29]), .o_cout(cout6[29]));
pu pu6_30 (.i_a(result5[29]), .i_b(~i_divisor[30]), .i_cin(cout6[29]), .i_carry_output(quotient[25]),
		.o_result(result6[30]), .o_cout(cout6[30]));
pu pu6_31 (.i_a(result5[30]), .i_b(~i_divisor[31]), .i_cin(cout6[30]), .i_carry_output(quotient[25]),
		.o_cout(quotient[25]));

// Row 7
pu pu7_0 (.i_a(i_dividend[24]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[24]),
         .o_result(result7[0]), .o_cout(cout7[0]));
pu pu7_1 (.i_a(result6[0]), .i_b(~i_divisor[1]), .i_cin(cout7[0]), .i_carry_output(quotient[24]),
		.o_result(result7[1]), .o_cout(cout7[1]));
pu pu7_2 (.i_a(result6[1]), .i_b(~i_divisor[2]), .i_cin(cout7[1]), .i_carry_output(quotient[24]),
		.o_result(result7[2]), .o_cout(cout7[2]));
pu pu7_3 (.i_a(result6[2]), .i_b(~i_divisor[3]), .i_cin(cout7[2]), .i_carry_output(quotient[24]),
		.o_result(result7[3]), .o_cout(cout7[3]));
pu pu7_4 (.i_a(result6[3]), .i_b(~i_divisor[4]), .i_cin(cout7[3]), .i_carry_output(quotient[24]),
		.o_result(result7[4]), .o_cout(cout7[4]));
pu pu7_5 (.i_a(result6[4]), .i_b(~i_divisor[5]), .i_cin(cout7[4]), .i_carry_output(quotient[24]),
		.o_result(result7[5]), .o_cout(cout7[5]));
pu pu7_6 (.i_a(result6[5]), .i_b(~i_divisor[6]), .i_cin(cout7[5]), .i_carry_output(quotient[24]),
		.o_result(result7[6]), .o_cout(cout7[6]));
pu pu7_7 (.i_a(result6[6]), .i_b(~i_divisor[7]), .i_cin(cout7[6]), .i_carry_output(quotient[24]),
		.o_result(result7[7]), .o_cout(cout7[7]));
pu pu7_8 (.i_a(result6[7]), .i_b(~i_divisor[8]), .i_cin(cout7[7]), .i_carry_output(quotient[24]),
		.o_result(result7[8]), .o_cout(cout7[8]));
pu pu7_9 (.i_a(result6[8]), .i_b(~i_divisor[9]), .i_cin(cout7[8]), .i_carry_output(quotient[24]),
		.o_result(result7[9]), .o_cout(cout7[9]));
pu pu7_10 (.i_a(result6[9]), .i_b(~i_divisor[10]), .i_cin(cout7[9]), .i_carry_output(quotient[24]),
		.o_result(result7[10]), .o_cout(cout7[10]));
pu pu7_11 (.i_a(result6[10]), .i_b(~i_divisor[11]), .i_cin(cout7[10]), .i_carry_output(quotient[24]),
		.o_result(result7[11]), .o_cout(cout7[11]));
pu pu7_12 (.i_a(result6[11]), .i_b(~i_divisor[12]), .i_cin(cout7[11]), .i_carry_output(quotient[24]),
		.o_result(result7[12]), .o_cout(cout7[12]));
pu pu7_13 (.i_a(result6[12]), .i_b(~i_divisor[13]), .i_cin(cout7[12]), .i_carry_output(quotient[24]),
		.o_result(result7[13]), .o_cout(cout7[13]));
pu pu7_14 (.i_a(result6[13]), .i_b(~i_divisor[14]), .i_cin(cout7[13]), .i_carry_output(quotient[24]),
		.o_result(result7[14]), .o_cout(cout7[14]));
pu pu7_15 (.i_a(result6[14]), .i_b(~i_divisor[15]), .i_cin(cout7[14]), .i_carry_output(quotient[24]),
		.o_result(result7[15]), .o_cout(cout7[15]));
pu pu7_16 (.i_a(result6[15]), .i_b(~i_divisor[16]), .i_cin(cout7[15]), .i_carry_output(quotient[24]),
		.o_result(result7[16]), .o_cout(cout7[16]));
pu pu7_17 (.i_a(result6[16]), .i_b(~i_divisor[17]), .i_cin(cout7[16]), .i_carry_output(quotient[24]),
		.o_result(result7[17]), .o_cout(cout7[17]));
pu pu7_18 (.i_a(result6[17]), .i_b(~i_divisor[18]), .i_cin(cout7[17]), .i_carry_output(quotient[24]),
		.o_result(result7[18]), .o_cout(cout7[18]));
pu pu7_19 (.i_a(result6[18]), .i_b(~i_divisor[19]), .i_cin(cout7[18]), .i_carry_output(quotient[24]),
		.o_result(result7[19]), .o_cout(cout7[19]));
pu pu7_20 (.i_a(result6[19]), .i_b(~i_divisor[20]), .i_cin(cout7[19]), .i_carry_output(quotient[24]),
		.o_result(result7[20]), .o_cout(cout7[20]));
pu pu7_21 (.i_a(result6[20]), .i_b(~i_divisor[21]), .i_cin(cout7[20]), .i_carry_output(quotient[24]),
		.o_result(result7[21]), .o_cout(cout7[21]));
pu pu7_22 (.i_a(result6[21]), .i_b(~i_divisor[22]), .i_cin(cout7[21]), .i_carry_output(quotient[24]),
		.o_result(result7[22]), .o_cout(cout7[22]));
pu pu7_23 (.i_a(result6[22]), .i_b(~i_divisor[23]), .i_cin(cout7[22]), .i_carry_output(quotient[24]),
		.o_result(result7[23]), .o_cout(cout7[23]));
pu pu7_24 (.i_a(result6[23]), .i_b(~i_divisor[24]), .i_cin(cout7[23]), .i_carry_output(quotient[24]),
		.o_result(result7[24]), .o_cout(cout7[24]));
pu pu7_25 (.i_a(result6[24]), .i_b(~i_divisor[25]), .i_cin(cout7[24]), .i_carry_output(quotient[24]),
		.o_result(result7[25]), .o_cout(cout7[25]));
pu pu7_26 (.i_a(result6[25]), .i_b(~i_divisor[26]), .i_cin(cout7[25]), .i_carry_output(quotient[24]),
		.o_result(result7[26]), .o_cout(cout7[26]));
pu pu7_27 (.i_a(result6[26]), .i_b(~i_divisor[27]), .i_cin(cout7[26]), .i_carry_output(quotient[24]),
		.o_result(result7[27]), .o_cout(cout7[27]));
pu pu7_28 (.i_a(result6[27]), .i_b(~i_divisor[28]), .i_cin(cout7[27]), .i_carry_output(quotient[24]),
		.o_result(result7[28]), .o_cout(cout7[28]));
pu pu7_29 (.i_a(result6[28]), .i_b(~i_divisor[29]), .i_cin(cout7[28]), .i_carry_output(quotient[24]),
		.o_result(result7[29]), .o_cout(cout7[29]));
pu pu7_30 (.i_a(result6[29]), .i_b(~i_divisor[30]), .i_cin(cout7[29]), .i_carry_output(quotient[24]),
		.o_result(result7[30]), .o_cout(cout7[30]));
pu pu7_31 (.i_a(result6[30]), .i_b(~i_divisor[31]), .i_cin(cout7[30]), .i_carry_output(quotient[24]),
		.o_cout(quotient[24]));

// Row 8
pu pu8_0 (.i_a(i_dividend[23]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[23]),
         .o_result(result8[0]), .o_cout(cout8[0]));
pu pu8_1 (.i_a(result7[0]), .i_b(~i_divisor[1]), .i_cin(cout8[0]), .i_carry_output(quotient[23]),
		.o_result(result8[1]), .o_cout(cout8[1]));
pu pu8_2 (.i_a(result7[1]), .i_b(~i_divisor[2]), .i_cin(cout8[1]), .i_carry_output(quotient[23]),
		.o_result(result8[2]), .o_cout(cout8[2]));
pu pu8_3 (.i_a(result7[2]), .i_b(~i_divisor[3]), .i_cin(cout8[2]), .i_carry_output(quotient[23]),
		.o_result(result8[3]), .o_cout(cout8[3]));
pu pu8_4 (.i_a(result7[3]), .i_b(~i_divisor[4]), .i_cin(cout8[3]), .i_carry_output(quotient[23]),
		.o_result(result8[4]), .o_cout(cout8[4]));
pu pu8_5 (.i_a(result7[4]), .i_b(~i_divisor[5]), .i_cin(cout8[4]), .i_carry_output(quotient[23]),
		.o_result(result8[5]), .o_cout(cout8[5]));
pu pu8_6 (.i_a(result7[5]), .i_b(~i_divisor[6]), .i_cin(cout8[5]), .i_carry_output(quotient[23]),
		.o_result(result8[6]), .o_cout(cout8[6]));
pu pu8_7 (.i_a(result7[6]), .i_b(~i_divisor[7]), .i_cin(cout8[6]), .i_carry_output(quotient[23]),
		.o_result(result8[7]), .o_cout(cout8[7]));
pu pu8_8 (.i_a(result7[7]), .i_b(~i_divisor[8]), .i_cin(cout8[7]), .i_carry_output(quotient[23]),
		.o_result(result8[8]), .o_cout(cout8[8]));
pu pu8_9 (.i_a(result7[8]), .i_b(~i_divisor[9]), .i_cin(cout8[8]), .i_carry_output(quotient[23]),
		.o_result(result8[9]), .o_cout(cout8[9]));
pu pu8_10 (.i_a(result7[9]), .i_b(~i_divisor[10]), .i_cin(cout8[9]), .i_carry_output(quotient[23]),
		.o_result(result8[10]), .o_cout(cout8[10]));
pu pu8_11 (.i_a(result7[10]), .i_b(~i_divisor[11]), .i_cin(cout8[10]), .i_carry_output(quotient[23]),
		.o_result(result8[11]), .o_cout(cout8[11]));
pu pu8_12 (.i_a(result7[11]), .i_b(~i_divisor[12]), .i_cin(cout8[11]), .i_carry_output(quotient[23]),
		.o_result(result8[12]), .o_cout(cout8[12]));
pu pu8_13 (.i_a(result7[12]), .i_b(~i_divisor[13]), .i_cin(cout8[12]), .i_carry_output(quotient[23]),
		.o_result(result8[13]), .o_cout(cout8[13]));
pu pu8_14 (.i_a(result7[13]), .i_b(~i_divisor[14]), .i_cin(cout8[13]), .i_carry_output(quotient[23]),
		.o_result(result8[14]), .o_cout(cout8[14]));
pu pu8_15 (.i_a(result7[14]), .i_b(~i_divisor[15]), .i_cin(cout8[14]), .i_carry_output(quotient[23]),
		.o_result(result8[15]), .o_cout(cout8[15]));
pu pu8_16 (.i_a(result7[15]), .i_b(~i_divisor[16]), .i_cin(cout8[15]), .i_carry_output(quotient[23]),
		.o_result(result8[16]), .o_cout(cout8[16]));
pu pu8_17 (.i_a(result7[16]), .i_b(~i_divisor[17]), .i_cin(cout8[16]), .i_carry_output(quotient[23]),
		.o_result(result8[17]), .o_cout(cout8[17]));
pu pu8_18 (.i_a(result7[17]), .i_b(~i_divisor[18]), .i_cin(cout8[17]), .i_carry_output(quotient[23]),
		.o_result(result8[18]), .o_cout(cout8[18]));
pu pu8_19 (.i_a(result7[18]), .i_b(~i_divisor[19]), .i_cin(cout8[18]), .i_carry_output(quotient[23]),
		.o_result(result8[19]), .o_cout(cout8[19]));
pu pu8_20 (.i_a(result7[19]), .i_b(~i_divisor[20]), .i_cin(cout8[19]), .i_carry_output(quotient[23]),
		.o_result(result8[20]), .o_cout(cout8[20]));
pu pu8_21 (.i_a(result7[20]), .i_b(~i_divisor[21]), .i_cin(cout8[20]), .i_carry_output(quotient[23]),
		.o_result(result8[21]), .o_cout(cout8[21]));
pu pu8_22 (.i_a(result7[21]), .i_b(~i_divisor[22]), .i_cin(cout8[21]), .i_carry_output(quotient[23]),
		.o_result(result8[22]), .o_cout(cout8[22]));
pu pu8_23 (.i_a(result7[22]), .i_b(~i_divisor[23]), .i_cin(cout8[22]), .i_carry_output(quotient[23]),
		.o_result(result8[23]), .o_cout(cout8[23]));
pu pu8_24 (.i_a(result7[23]), .i_b(~i_divisor[24]), .i_cin(cout8[23]), .i_carry_output(quotient[23]),
		.o_result(result8[24]), .o_cout(cout8[24]));
pu pu8_25 (.i_a(result7[24]), .i_b(~i_divisor[25]), .i_cin(cout8[24]), .i_carry_output(quotient[23]),
		.o_result(result8[25]), .o_cout(cout8[25]));
pu pu8_26 (.i_a(result7[25]), .i_b(~i_divisor[26]), .i_cin(cout8[25]), .i_carry_output(quotient[23]),
		.o_result(result8[26]), .o_cout(cout8[26]));
pu pu8_27 (.i_a(result7[26]), .i_b(~i_divisor[27]), .i_cin(cout8[26]), .i_carry_output(quotient[23]),
		.o_result(result8[27]), .o_cout(cout8[27]));
pu pu8_28 (.i_a(result7[27]), .i_b(~i_divisor[28]), .i_cin(cout8[27]), .i_carry_output(quotient[23]),
		.o_result(result8[28]), .o_cout(cout8[28]));
pu pu8_29 (.i_a(result7[28]), .i_b(~i_divisor[29]), .i_cin(cout8[28]), .i_carry_output(quotient[23]),
		.o_result(result8[29]), .o_cout(cout8[29]));
pu pu8_30 (.i_a(result7[29]), .i_b(~i_divisor[30]), .i_cin(cout8[29]), .i_carry_output(quotient[23]),
		.o_result(result8[30]), .o_cout(cout8[30]));
pu pu8_31 (.i_a(result7[30]), .i_b(~i_divisor[31]), .i_cin(cout8[30]), .i_carry_output(quotient[23]),
		.o_cout(quotient[23]));

// Row 9
pu pu9_0 (.i_a(i_dividend[22]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[22]),
         .o_result(result9[0]), .o_cout(cout9[0]));
pu pu91 (.i_a(result8[0]), .i_b(~i_divisor[1]), .i_cin(cout9[0]), .i_carry_output(quotient[22]),
		.o_result(result9[1]), .o_cout(cout9[1]));
pu pu9_2 (.i_a(result8[1]), .i_b(~i_divisor[2]), .i_cin(cout9[1]), .i_carry_output(quotient[22]),
		.o_result(result9[2]), .o_cout(cout9[2]));
pu pu9_3 (.i_a(result8[2]), .i_b(~i_divisor[3]), .i_cin(cout9[2]), .i_carry_output(quotient[22]),
		.o_result(result9[3]), .o_cout(cout9[3]));
pu pu9_4 (.i_a(result8[3]), .i_b(~i_divisor[4]), .i_cin(cout9[3]), .i_carry_output(quotient[22]),
		.o_result(result9[4]), .o_cout(cout9[4]));
pu pu9_5 (.i_a(result8[4]), .i_b(~i_divisor[5]), .i_cin(cout9[4]), .i_carry_output(quotient[22]),
		.o_result(result9[5]), .o_cout(cout9[5]));
pu pu9_6 (.i_a(result8[5]), .i_b(~i_divisor[6]), .i_cin(cout9[5]), .i_carry_output(quotient[22]),
		.o_result(result9[6]), .o_cout(cout9[6]));
pu pu9_7 (.i_a(result8[6]), .i_b(~i_divisor[7]), .i_cin(cout9[6]), .i_carry_output(quotient[22]),
		.o_result(result9[7]), .o_cout(cout9[7]));
pu pu9_8 (.i_a(result8[7]), .i_b(~i_divisor[8]), .i_cin(cout9[7]), .i_carry_output(quotient[22]),
		.o_result(result9[8]), .o_cout(cout9[8]));
pu pu9_9 (.i_a(result8[8]), .i_b(~i_divisor[9]), .i_cin(cout9[8]), .i_carry_output(quotient[22]),
		.o_result(result9[9]), .o_cout(cout9[9]));
pu pu9_10 (.i_a(result8[9]), .i_b(~i_divisor[10]), .i_cin(cout9[9]), .i_carry_output(quotient[22]),
		.o_result(result9[10]), .o_cout(cout9[10]));
pu pu9_11 (.i_a(result8[10]), .i_b(~i_divisor[11]), .i_cin(cout9[10]), .i_carry_output(quotient[22]),
		.o_result(result9[11]), .o_cout(cout9[11]));
pu pu9_12 (.i_a(result8[11]), .i_b(~i_divisor[12]), .i_cin(cout9[11]), .i_carry_output(quotient[22]),
		.o_result(result9[12]), .o_cout(cout9[12]));
pu pu9_13 (.i_a(result8[12]), .i_b(~i_divisor[13]), .i_cin(cout9[12]), .i_carry_output(quotient[22]),
		.o_result(result9[13]), .o_cout(cout9[13]));
pu pu9_14 (.i_a(result8[13]), .i_b(~i_divisor[14]), .i_cin(cout9[13]), .i_carry_output(quotient[22]),
		.o_result(result9[14]), .o_cout(cout9[14]));
pu pu9_15 (.i_a(result8[14]), .i_b(~i_divisor[15]), .i_cin(cout9[14]), .i_carry_output(quotient[22]),
		.o_result(result9[15]), .o_cout(cout9[15]));
pu pu9_16 (.i_a(result8[15]), .i_b(~i_divisor[16]), .i_cin(cout9[15]), .i_carry_output(quotient[22]),
		.o_result(result9[16]), .o_cout(cout9[16]));
pu pu9_17 (.i_a(result8[16]), .i_b(~i_divisor[17]), .i_cin(cout9[16]), .i_carry_output(quotient[22]),
		.o_result(result9[17]), .o_cout(cout9[17]));
pu pu9_18 (.i_a(result8[17]), .i_b(~i_divisor[18]), .i_cin(cout9[17]), .i_carry_output(quotient[22]),
		.o_result(result9[18]), .o_cout(cout9[18]));
pu pu9_19 (.i_a(result8[18]), .i_b(~i_divisor[19]), .i_cin(cout9[18]), .i_carry_output(quotient[22]),
		.o_result(result9[19]), .o_cout(cout9[19]));
pu pu9_20 (.i_a(result8[19]), .i_b(~i_divisor[20]), .i_cin(cout9[19]), .i_carry_output(quotient[22]),
		.o_result(result9[20]), .o_cout(cout9[20]));
pu pu9_21 (.i_a(result8[20]), .i_b(~i_divisor[21]), .i_cin(cout9[20]), .i_carry_output(quotient[22]),
		.o_result(result9[21]), .o_cout(cout9[21]));
pu pu9_22 (.i_a(result8[21]), .i_b(~i_divisor[22]), .i_cin(cout9[21]), .i_carry_output(quotient[22]),
		.o_result(result9[22]), .o_cout(cout9[22]));
pu pu9_23 (.i_a(result8[22]), .i_b(~i_divisor[23]), .i_cin(cout9[22]), .i_carry_output(quotient[22]),
		.o_result(result9[23]), .o_cout(cout9[23]));
pu pu9_24 (.i_a(result8[23]), .i_b(~i_divisor[24]), .i_cin(cout9[23]), .i_carry_output(quotient[22]),
		.o_result(result9[24]), .o_cout(cout9[24]));
pu pu9_25 (.i_a(result8[24]), .i_b(~i_divisor[25]), .i_cin(cout9[24]), .i_carry_output(quotient[22]),
		.o_result(result9[25]), .o_cout(cout9[25]));
pu pu9_26 (.i_a(result8[25]), .i_b(~i_divisor[26]), .i_cin(cout9[25]), .i_carry_output(quotient[22]),
		.o_result(result9[26]), .o_cout(cout9[26]));
pu pu9_27 (.i_a(result8[26]), .i_b(~i_divisor[27]), .i_cin(cout9[26]), .i_carry_output(quotient[22]),
		.o_result(result9[27]), .o_cout(cout9[27]));
pu pu9_28 (.i_a(result8[27]), .i_b(~i_divisor[28]), .i_cin(cout9[27]), .i_carry_output(quotient[22]),
		.o_result(result9[28]), .o_cout(cout9[28]));
pu pu9_29 (.i_a(result8[28]), .i_b(~i_divisor[29]), .i_cin(cout9[28]), .i_carry_output(quotient[22]),
		.o_result(result9[29]), .o_cout(cout9[29]));
pu pu9_30 (.i_a(result8[29]), .i_b(~i_divisor[30]), .i_cin(cout9[29]), .i_carry_output(quotient[22]),
		.o_result(result9[30]), .o_cout(cout9[30]));
pu pu9_31 (.i_a(result8[30]), .i_b(~i_divisor[31]), .i_cin(cout9[30]), .i_carry_output(quotient[22]),
		.o_cout(quotient[22]));

// Row 10
pu pu100 (.i_a(i_dividend[21]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[21]),
         .o_result(result10[0]), .o_cout(cout10[0]));
pu pu10_1 (.i_a(result9[0]), .i_b(~i_divisor[1]), .i_cin(cout10[0]), .i_carry_output(quotient[21]),
		.o_result(result10[1]), .o_cout(cout10[1]));
pu pu10_2 (.i_a(result9[1]), .i_b(~i_divisor[2]), .i_cin(cout10[1]), .i_carry_output(quotient[21]),
		.o_result(result10[2]), .o_cout(cout10[2]));
pu pu10_3 (.i_a(result9[2]), .i_b(~i_divisor[3]), .i_cin(cout10[2]), .i_carry_output(quotient[21]),
		.o_result(result10[3]), .o_cout(cout10[3]));
pu pu10_4 (.i_a(result9[3]), .i_b(~i_divisor[4]), .i_cin(cout10[3]), .i_carry_output(quotient[21]),
		.o_result(result10[4]), .o_cout(cout10[4]));
pu pu10_5 (.i_a(result9[4]), .i_b(~i_divisor[5]), .i_cin(cout10[4]), .i_carry_output(quotient[21]),
		.o_result(result10[5]), .o_cout(cout10[5]));
pu pu10_6 (.i_a(result9[5]), .i_b(~i_divisor[6]), .i_cin(cout10[5]), .i_carry_output(quotient[21]),
		.o_result(result10[6]), .o_cout(cout10[6]));
pu pu10_7 (.i_a(result9[6]), .i_b(~i_divisor[7]), .i_cin(cout10[6]), .i_carry_output(quotient[21]),
		.o_result(result10[7]), .o_cout(cout10[7]));
pu pu10_8 (.i_a(result9[7]), .i_b(~i_divisor[8]), .i_cin(cout10[7]), .i_carry_output(quotient[21]),
		.o_result(result10[8]), .o_cout(cout10[8]));
pu pu10_9 (.i_a(result9[8]), .i_b(~i_divisor[9]), .i_cin(cout10[8]), .i_carry_output(quotient[21]),
		.o_result(result10[9]), .o_cout(cout10[9]));
pu pu10_10 (.i_a(result9[9]), .i_b(~i_divisor[10]), .i_cin(cout10[9]), .i_carry_output(quotient[21]),
		.o_result(result10[10]), .o_cout(cout10[10]));
pu pu10_11 (.i_a(result9[10]), .i_b(~i_divisor[11]), .i_cin(cout10[10]), .i_carry_output(quotient[21]),
		.o_result(result10[11]), .o_cout(cout10[11]));
pu pu10_12 (.i_a(result9[11]), .i_b(~i_divisor[12]), .i_cin(cout10[11]), .i_carry_output(quotient[21]),
		.o_result(result10[12]), .o_cout(cout10[12]));
pu pu10_13 (.i_a(result9[12]), .i_b(~i_divisor[13]), .i_cin(cout10[12]), .i_carry_output(quotient[21]),
		.o_result(result10[13]), .o_cout(cout10[13]));
pu pu10_14 (.i_a(result9[13]), .i_b(~i_divisor[14]), .i_cin(cout10[13]), .i_carry_output(quotient[21]),
		.o_result(result10[14]), .o_cout(cout10[14]));
pu pu10_15 (.i_a(result9[14]), .i_b(~i_divisor[15]), .i_cin(cout10[14]), .i_carry_output(quotient[21]),
		.o_result(result10[15]), .o_cout(cout10[15]));
pu pu10_16 (.i_a(result9[15]), .i_b(~i_divisor[16]), .i_cin(cout10[15]), .i_carry_output(quotient[21]),
		.o_result(result10[16]), .o_cout(cout10[16]));
pu pu10_17 (.i_a(result9[16]), .i_b(~i_divisor[17]), .i_cin(cout10[16]), .i_carry_output(quotient[21]),
		.o_result(result10[17]), .o_cout(cout10[17]));
pu pu10_18 (.i_a(result9[17]), .i_b(~i_divisor[18]), .i_cin(cout10[17]), .i_carry_output(quotient[21]),
		.o_result(result10[18]), .o_cout(cout10[18]));
pu pu10_19 (.i_a(result9[18]), .i_b(~i_divisor[19]), .i_cin(cout10[18]), .i_carry_output(quotient[21]),
		.o_result(result10[19]), .o_cout(cout10[19]));
pu pu10_20 (.i_a(result9[19]), .i_b(~i_divisor[20]), .i_cin(cout10[19]), .i_carry_output(quotient[21]),
		.o_result(result10[20]), .o_cout(cout10[20]));
pu pu10_21 (.i_a(result9[20]), .i_b(~i_divisor[21]), .i_cin(cout10[20]), .i_carry_output(quotient[21]),
		.o_result(result10[21]), .o_cout(cout10[21]));
pu pu10_22 (.i_a(result9[21]), .i_b(~i_divisor[22]), .i_cin(cout10[21]), .i_carry_output(quotient[21]),
		.o_result(result10[22]), .o_cout(cout10[22]));
pu pu10_23 (.i_a(result9[22]), .i_b(~i_divisor[23]), .i_cin(cout10[22]), .i_carry_output(quotient[21]),
		.o_result(result10[23]), .o_cout(cout10[23]));
pu pu10_24 (.i_a(result9[23]), .i_b(~i_divisor[24]), .i_cin(cout10[23]), .i_carry_output(quotient[21]),
		.o_result(result10[24]), .o_cout(cout10[24]));
pu pu10_25 (.i_a(result9[24]), .i_b(~i_divisor[25]), .i_cin(cout10[24]), .i_carry_output(quotient[21]),
		.o_result(result10[25]), .o_cout(cout10[25]));
pu pu10_26 (.i_a(result9[25]), .i_b(~i_divisor[26]), .i_cin(cout10[25]), .i_carry_output(quotient[21]),
		.o_result(result10[26]), .o_cout(cout10[26]));
pu pu10_27 (.i_a(result9[26]), .i_b(~i_divisor[27]), .i_cin(cout10[26]), .i_carry_output(quotient[21]),
		.o_result(result10[27]), .o_cout(cout10[27]));
pu pu10_28 (.i_a(result9[27]), .i_b(~i_divisor[28]), .i_cin(cout10[27]), .i_carry_output(quotient[21]),
		.o_result(result10[28]), .o_cout(cout10[28]));
pu pu10_29 (.i_a(result9[28]), .i_b(~i_divisor[29]), .i_cin(cout10[28]), .i_carry_output(quotient[21]),
		.o_result(result10[29]), .o_cout(cout10[29]));
pu pu10_30 (.i_a(result9[29]), .i_b(~i_divisor[30]), .i_cin(cout10[29]), .i_carry_output(quotient[21]),
		.o_result(result10[30]), .o_cout(cout10[30]));
pu pu10_31 (.i_a(result9[30]), .i_b(~i_divisor[31]), .i_cin(cout10[30]), .i_carry_output(quotient[21]),
		.o_cout(quotient[21]));

// Row 11
pu pu11_0 (.i_a(i_dividend[20]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[20]),
         .o_result(result11[0]), .o_cout(cout11[0]));
pu pu11_1 (.i_a(result10[0]), .i_b(~i_divisor[1]), .i_cin(cout11[0]), .i_carry_output(quotient[20]),
		.o_result(result11[1]), .o_cout(cout11[1]));
pu pu11_2 (.i_a(result10[1]), .i_b(~i_divisor[2]), .i_cin(cout11[1]), .i_carry_output(quotient[20]),
		.o_result(result11[2]), .o_cout(cout11[2]));
pu pu11_3 (.i_a(result10[2]), .i_b(~i_divisor[3]), .i_cin(cout11[2]), .i_carry_output(quotient[20]),
		.o_result(result11[3]), .o_cout(cout11[3]));
pu pu11_4 (.i_a(result10[3]), .i_b(~i_divisor[4]), .i_cin(cout11[3]), .i_carry_output(quotient[20]),
		.o_result(result11[4]), .o_cout(cout11[4]));
pu pu11_5 (.i_a(result10[4]), .i_b(~i_divisor[5]), .i_cin(cout11[4]), .i_carry_output(quotient[20]),
		.o_result(result11[5]), .o_cout(cout11[5]));
pu pu11_6 (.i_a(result10[5]), .i_b(~i_divisor[6]), .i_cin(cout11[5]), .i_carry_output(quotient[20]),
		.o_result(result11[6]), .o_cout(cout11[6]));
pu pu11_7 (.i_a(result10[6]), .i_b(~i_divisor[7]), .i_cin(cout11[6]), .i_carry_output(quotient[20]),
		.o_result(result11[7]), .o_cout(cout11[7]));
pu pu11_8 (.i_a(result10[7]), .i_b(~i_divisor[8]), .i_cin(cout11[7]), .i_carry_output(quotient[20]),
		.o_result(result11[8]), .o_cout(cout11[8]));
pu pu11_9 (.i_a(result10[8]), .i_b(~i_divisor[9]), .i_cin(cout11[8]), .i_carry_output(quotient[20]),
		.o_result(result11[9]), .o_cout(cout11[9]));
pu pu11_10 (.i_a(result10[9]), .i_b(~i_divisor[10]), .i_cin(cout11[9]), .i_carry_output(quotient[20]),
		.o_result(result11[10]), .o_cout(cout11[10]));
pu pu11_11 (.i_a(result10[10]), .i_b(~i_divisor[11]), .i_cin(cout11[10]), .i_carry_output(quotient[20]),
		.o_result(result11[11]), .o_cout(cout11[11]));
pu pu11_12 (.i_a(result10[11]), .i_b(~i_divisor[12]), .i_cin(cout11[11]), .i_carry_output(quotient[20]),
		.o_result(result11[12]), .o_cout(cout11[12]));
pu pu11_13 (.i_a(result10[12]), .i_b(~i_divisor[13]), .i_cin(cout11[12]), .i_carry_output(quotient[20]),
		.o_result(result11[13]), .o_cout(cout11[13]));
pu pu11_14 (.i_a(result10[13]), .i_b(~i_divisor[14]), .i_cin(cout11[13]), .i_carry_output(quotient[20]),
		.o_result(result11[14]), .o_cout(cout11[14]));
pu pu11_15 (.i_a(result10[14]), .i_b(~i_divisor[15]), .i_cin(cout11[14]), .i_carry_output(quotient[20]),
		.o_result(result11[15]), .o_cout(cout11[15]));
pu pu11_16 (.i_a(result10[15]), .i_b(~i_divisor[16]), .i_cin(cout11[15]), .i_carry_output(quotient[20]),
		.o_result(result11[16]), .o_cout(cout11[16]));
pu pu11_17 (.i_a(result10[16]), .i_b(~i_divisor[17]), .i_cin(cout11[16]), .i_carry_output(quotient[20]),
		.o_result(result11[17]), .o_cout(cout11[17]));
pu pu11_18 (.i_a(result10[17]), .i_b(~i_divisor[18]), .i_cin(cout11[17]), .i_carry_output(quotient[20]),
		.o_result(result11[18]), .o_cout(cout11[18]));
pu pu11_19 (.i_a(result10[18]), .i_b(~i_divisor[19]), .i_cin(cout11[18]), .i_carry_output(quotient[20]),
		.o_result(result11[19]), .o_cout(cout11[19]));
pu pu11_20 (.i_a(result10[19]), .i_b(~i_divisor[20]), .i_cin(cout11[19]), .i_carry_output(quotient[20]),
		.o_result(result11[20]), .o_cout(cout11[20]));
pu pu11_21 (.i_a(result10[20]), .i_b(~i_divisor[21]), .i_cin(cout11[20]), .i_carry_output(quotient[20]),
		.o_result(result11[21]), .o_cout(cout11[21]));
pu pu11_22 (.i_a(result10[21]), .i_b(~i_divisor[22]), .i_cin(cout11[21]), .i_carry_output(quotient[20]),
		.o_result(result11[22]), .o_cout(cout11[22]));
pu pu11_23 (.i_a(result10[22]), .i_b(~i_divisor[23]), .i_cin(cout11[22]), .i_carry_output(quotient[20]),
		.o_result(result11[23]), .o_cout(cout11[23]));
pu pu11_24 (.i_a(result10[23]), .i_b(~i_divisor[24]), .i_cin(cout11[23]), .i_carry_output(quotient[20]),
		.o_result(result11[24]), .o_cout(cout11[24]));
pu pu11_25 (.i_a(result10[24]), .i_b(~i_divisor[25]), .i_cin(cout11[24]), .i_carry_output(quotient[20]),
		.o_result(result11[25]), .o_cout(cout11[25]));
pu pu11_26 (.i_a(result10[25]), .i_b(~i_divisor[26]), .i_cin(cout11[25]), .i_carry_output(quotient[20]),
		.o_result(result11[26]), .o_cout(cout11[26]));
pu pu11_27 (.i_a(result10[26]), .i_b(~i_divisor[27]), .i_cin(cout11[26]), .i_carry_output(quotient[20]),
		.o_result(result11[27]), .o_cout(cout11[27]));
pu pu11_28 (.i_a(result10[27]), .i_b(~i_divisor[28]), .i_cin(cout11[27]), .i_carry_output(quotient[20]),
		.o_result(result11[28]), .o_cout(cout11[28]));
pu pu11_29 (.i_a(result10[28]), .i_b(~i_divisor[29]), .i_cin(cout11[28]), .i_carry_output(quotient[20]),
		.o_result(result11[29]), .o_cout(cout11[29]));
pu pu11_30 (.i_a(result10[29]), .i_b(~i_divisor[30]), .i_cin(cout11[29]), .i_carry_output(quotient[20]),
		.o_result(result11[30]), .o_cout(cout11[30]));
pu pu11_31 (.i_a(result10[30]), .i_b(~i_divisor[31]), .i_cin(cout11[30]), .i_carry_output(quotient[20]),
		.o_cout(quotient[20]));

// Row 12
pu pu12_0 (.i_a(i_dividend[19]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[19]),
         .o_result(result12[0]), .o_cout(cout12[0]));
pu pu12_1 (.i_a(result11[0]), .i_b(~i_divisor[1]), .i_cin(cout12[0]), .i_carry_output(quotient[19]),
		.o_result(result12[1]), .o_cout(cout12[1]));
pu pu12_2 (.i_a(result11[1]), .i_b(~i_divisor[2]), .i_cin(cout12[1]), .i_carry_output(quotient[19]),
		.o_result(result12[2]), .o_cout(cout12[2]));
pu pu12_3 (.i_a(result11[2]), .i_b(~i_divisor[3]), .i_cin(cout12[2]), .i_carry_output(quotient[19]),
		.o_result(result12[3]), .o_cout(cout12[3]));
pu pu12_4 (.i_a(result11[3]), .i_b(~i_divisor[4]), .i_cin(cout12[3]), .i_carry_output(quotient[19]),
		.o_result(result12[4]), .o_cout(cout12[4]));
pu pu12_5 (.i_a(result11[4]), .i_b(~i_divisor[5]), .i_cin(cout12[4]), .i_carry_output(quotient[19]),
		.o_result(result12[5]), .o_cout(cout12[5]));
pu pu12_6 (.i_a(result11[5]), .i_b(~i_divisor[6]), .i_cin(cout12[5]), .i_carry_output(quotient[19]),
		.o_result(result12[6]), .o_cout(cout12[6]));
pu pu12_7 (.i_a(result11[6]), .i_b(~i_divisor[7]), .i_cin(cout12[6]), .i_carry_output(quotient[19]),
		.o_result(result12[7]), .o_cout(cout12[7]));
pu pu12_8 (.i_a(result11[7]), .i_b(~i_divisor[8]), .i_cin(cout12[7]), .i_carry_output(quotient[19]),
		.o_result(result12[8]), .o_cout(cout12[8]));
pu pu12_9 (.i_a(result11[8]), .i_b(~i_divisor[9]), .i_cin(cout12[8]), .i_carry_output(quotient[19]),
		.o_result(result12[9]), .o_cout(cout12[9]));
pu pu12_10 (.i_a(result11[9]), .i_b(~i_divisor[10]), .i_cin(cout12[9]), .i_carry_output(quotient[19]),
		.o_result(result12[10]), .o_cout(cout12[10]));
pu pu12_11 (.i_a(result11[10]), .i_b(~i_divisor[11]), .i_cin(cout12[10]), .i_carry_output(quotient[19]),
		.o_result(result12[11]), .o_cout(cout12[11]));
pu pu12_12 (.i_a(result11[11]), .i_b(~i_divisor[12]), .i_cin(cout12[11]), .i_carry_output(quotient[19]),
		.o_result(result12[12]), .o_cout(cout12[12]));
pu pu12_13 (.i_a(result11[12]), .i_b(~i_divisor[13]), .i_cin(cout12[12]), .i_carry_output(quotient[19]),
		.o_result(result12[13]), .o_cout(cout12[13]));
pu pu12_14 (.i_a(result11[13]), .i_b(~i_divisor[14]), .i_cin(cout12[13]), .i_carry_output(quotient[19]),
		.o_result(result12[14]), .o_cout(cout12[14]));
pu pu12_15 (.i_a(result11[14]), .i_b(~i_divisor[15]), .i_cin(cout12[14]), .i_carry_output(quotient[19]),
		.o_result(result12[15]), .o_cout(cout12[15]));
pu pu12_16 (.i_a(result11[15]), .i_b(~i_divisor[16]), .i_cin(cout12[15]), .i_carry_output(quotient[19]),
		.o_result(result12[16]), .o_cout(cout12[16]));
pu pu12_17 (.i_a(result11[16]), .i_b(~i_divisor[17]), .i_cin(cout12[16]), .i_carry_output(quotient[19]),
		.o_result(result12[17]), .o_cout(cout12[17]));
pu pu12_18 (.i_a(result11[17]), .i_b(~i_divisor[18]), .i_cin(cout12[17]), .i_carry_output(quotient[19]),
		.o_result(result12[18]), .o_cout(cout12[18]));
pu pu12_19 (.i_a(result11[18]), .i_b(~i_divisor[19]), .i_cin(cout12[18]), .i_carry_output(quotient[19]),
		.o_result(result12[19]), .o_cout(cout12[19]));
pu pu12_20 (.i_a(result11[19]), .i_b(~i_divisor[20]), .i_cin(cout12[19]), .i_carry_output(quotient[19]),
		.o_result(result12[20]), .o_cout(cout12[20]));
pu pu12_21 (.i_a(result11[20]), .i_b(~i_divisor[21]), .i_cin(cout12[20]), .i_carry_output(quotient[19]),
		.o_result(result12[21]), .o_cout(cout12[21]));
pu pu12_22 (.i_a(result11[21]), .i_b(~i_divisor[22]), .i_cin(cout12[21]), .i_carry_output(quotient[19]),
		.o_result(result12[22]), .o_cout(cout12[22]));
pu pu12_23 (.i_a(result11[22]), .i_b(~i_divisor[23]), .i_cin(cout12[22]), .i_carry_output(quotient[19]),
		.o_result(result12[23]), .o_cout(cout12[23]));
pu pu12_24 (.i_a(result11[23]), .i_b(~i_divisor[24]), .i_cin(cout12[23]), .i_carry_output(quotient[19]),
		.o_result(result12[24]), .o_cout(cout12[24]));
pu pu12_25 (.i_a(result11[24]), .i_b(~i_divisor[25]), .i_cin(cout12[24]), .i_carry_output(quotient[19]),
		.o_result(result12[25]), .o_cout(cout12[25]));
pu pu12_26 (.i_a(result11[25]), .i_b(~i_divisor[26]), .i_cin(cout12[25]), .i_carry_output(quotient[19]),
		.o_result(result12[26]), .o_cout(cout12[26]));
pu pu12_27 (.i_a(result11[26]), .i_b(~i_divisor[27]), .i_cin(cout12[26]), .i_carry_output(quotient[19]),
		.o_result(result12[27]), .o_cout(cout12[27]));
pu pu12_28 (.i_a(result11[27]), .i_b(~i_divisor[28]), .i_cin(cout12[27]), .i_carry_output(quotient[19]),
		.o_result(result12[28]), .o_cout(cout12[28]));
pu pu12_29 (.i_a(result11[28]), .i_b(~i_divisor[29]), .i_cin(cout12[28]), .i_carry_output(quotient[19]),
		.o_result(result12[29]), .o_cout(cout12[29]));
pu pu12_30 (.i_a(result11[29]), .i_b(~i_divisor[30]), .i_cin(cout12[29]), .i_carry_output(quotient[19]),
		.o_result(result12[30]), .o_cout(cout12[30]));
pu pu12_31 (.i_a(result11[30]), .i_b(~i_divisor[31]), .i_cin(cout12[30]), .i_carry_output(quotient[19]),
		.o_cout(quotient[19]));

// Row 13
pu pu13_0 (.i_a(i_dividend[18]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[18]),
         .o_result(result13[0]), .o_cout(cout13[0]));
pu pu13_1 (.i_a(result12[0]), .i_b(~i_divisor[1]), .i_cin(cout13[0]), .i_carry_output(quotient[18]),
		.o_result(result13[1]), .o_cout(cout13[1]));
pu pu13_2 (.i_a(result12[1]), .i_b(~i_divisor[2]), .i_cin(cout13[1]), .i_carry_output(quotient[18]),
		.o_result(result13[2]), .o_cout(cout13[2]));
pu pu13_3 (.i_a(result12[2]), .i_b(~i_divisor[3]), .i_cin(cout13[2]), .i_carry_output(quotient[18]),
		.o_result(result13[3]), .o_cout(cout13[3]));
pu pu13_4 (.i_a(result12[3]), .i_b(~i_divisor[4]), .i_cin(cout13[3]), .i_carry_output(quotient[18]),
		.o_result(result13[4]), .o_cout(cout13[4]));
pu pu13_5 (.i_a(result12[4]), .i_b(~i_divisor[5]), .i_cin(cout13[4]), .i_carry_output(quotient[18]),
		.o_result(result13[5]), .o_cout(cout13[5]));
pu pu13_6 (.i_a(result12[5]), .i_b(~i_divisor[6]), .i_cin(cout13[5]), .i_carry_output(quotient[18]),
		.o_result(result13[6]), .o_cout(cout13[6]));
pu pu13_7 (.i_a(result12[6]), .i_b(~i_divisor[7]), .i_cin(cout13[6]), .i_carry_output(quotient[18]),
		.o_result(result13[7]), .o_cout(cout13[7]));
pu pu13_8 (.i_a(result12[7]), .i_b(~i_divisor[8]), .i_cin(cout13[7]), .i_carry_output(quotient[18]),
		.o_result(result13[8]), .o_cout(cout13[8]));
pu pu13_9 (.i_a(result12[8]), .i_b(~i_divisor[9]), .i_cin(cout13[8]), .i_carry_output(quotient[18]),
		.o_result(result13[9]), .o_cout(cout13[9]));
pu pu13_10 (.i_a(result12[9]), .i_b(~i_divisor[10]), .i_cin(cout13[9]), .i_carry_output(quotient[18]),
		.o_result(result13[10]), .o_cout(cout13[10]));
pu pu13_11 (.i_a(result12[10]), .i_b(~i_divisor[11]), .i_cin(cout13[10]), .i_carry_output(quotient[18]),
		.o_result(result13[11]), .o_cout(cout13[11]));
pu pu13_12 (.i_a(result12[11]), .i_b(~i_divisor[12]), .i_cin(cout13[11]), .i_carry_output(quotient[18]),
		.o_result(result13[12]), .o_cout(cout13[12]));
pu pu13_13 (.i_a(result12[12]), .i_b(~i_divisor[13]), .i_cin(cout13[12]), .i_carry_output(quotient[18]),
		.o_result(result13[13]), .o_cout(cout13[13]));
pu pu13_14 (.i_a(result12[13]), .i_b(~i_divisor[14]), .i_cin(cout13[13]), .i_carry_output(quotient[18]),
		.o_result(result13[14]), .o_cout(cout13[14]));
pu pu13_15 (.i_a(result12[14]), .i_b(~i_divisor[15]), .i_cin(cout13[14]), .i_carry_output(quotient[18]),
		.o_result(result13[15]), .o_cout(cout13[15]));
pu pu13_16 (.i_a(result12[15]), .i_b(~i_divisor[16]), .i_cin(cout13[15]), .i_carry_output(quotient[18]),
		.o_result(result13[16]), .o_cout(cout13[16]));
pu pu13_17 (.i_a(result12[16]), .i_b(~i_divisor[17]), .i_cin(cout13[16]), .i_carry_output(quotient[18]),
		.o_result(result13[17]), .o_cout(cout13[17]));
pu pu13_18 (.i_a(result12[17]), .i_b(~i_divisor[18]), .i_cin(cout13[17]), .i_carry_output(quotient[18]),
		.o_result(result13[18]), .o_cout(cout13[18]));
pu pu13_19 (.i_a(result12[18]), .i_b(~i_divisor[19]), .i_cin(cout13[18]), .i_carry_output(quotient[18]),
		.o_result(result13[19]), .o_cout(cout13[19]));
pu pu13_20 (.i_a(result12[19]), .i_b(~i_divisor[20]), .i_cin(cout13[19]), .i_carry_output(quotient[18]),
		.o_result(result13[20]), .o_cout(cout13[20]));
pu pu13_21 (.i_a(result12[20]), .i_b(~i_divisor[21]), .i_cin(cout13[20]), .i_carry_output(quotient[18]),
		.o_result(result13[21]), .o_cout(cout13[21]));
pu pu13_22 (.i_a(result12[21]), .i_b(~i_divisor[22]), .i_cin(cout13[21]), .i_carry_output(quotient[18]),
		.o_result(result13[22]), .o_cout(cout13[22]));
pu pu13_23 (.i_a(result12[22]), .i_b(~i_divisor[23]), .i_cin(cout13[22]), .i_carry_output(quotient[18]),
		.o_result(result13[23]), .o_cout(cout13[23]));
pu pu13_24 (.i_a(result12[23]), .i_b(~i_divisor[24]), .i_cin(cout13[23]), .i_carry_output(quotient[18]),
		.o_result(result13[24]), .o_cout(cout13[24]));
pu pu13_25 (.i_a(result12[24]), .i_b(~i_divisor[25]), .i_cin(cout13[24]), .i_carry_output(quotient[18]),
		.o_result(result13[25]), .o_cout(cout13[25]));
pu pu13_26 (.i_a(result12[25]), .i_b(~i_divisor[26]), .i_cin(cout13[25]), .i_carry_output(quotient[18]),
		.o_result(result13[26]), .o_cout(cout13[26]));
pu pu13_27 (.i_a(result12[26]), .i_b(~i_divisor[27]), .i_cin(cout13[26]), .i_carry_output(quotient[18]),
		.o_result(result13[27]), .o_cout(cout13[27]));
pu pu13_28 (.i_a(result12[27]), .i_b(~i_divisor[28]), .i_cin(cout13[27]), .i_carry_output(quotient[18]),
		.o_result(result13[28]), .o_cout(cout13[28]));
pu pu13_29 (.i_a(result12[28]), .i_b(~i_divisor[29]), .i_cin(cout13[28]), .i_carry_output(quotient[18]),
		.o_result(result13[29]), .o_cout(cout13[29]));
pu pu13_30 (.i_a(result12[29]), .i_b(~i_divisor[30]), .i_cin(cout13[29]), .i_carry_output(quotient[18]),
		.o_result(result13[30]), .o_cout(cout13[30]));
pu pu13_31 (.i_a(result12[30]), .i_b(~i_divisor[31]), .i_cin(cout13[30]), .i_carry_output(quotient[18]),
		.o_cout(quotient[18]));

// Row 14
pu pu14_0 (.i_a(i_dividend[17]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[17]),
         .o_result(result14[0]), .o_cout(cout14[0]));
pu pu14_1 (.i_a(result13[0]), .i_b(~i_divisor[1]), .i_cin(cout14[0]), .i_carry_output(quotient[17]),
		.o_result(result14[1]), .o_cout(cout14[1]));
pu pu14_2 (.i_a(result13[1]), .i_b(~i_divisor[2]), .i_cin(cout14[1]), .i_carry_output(quotient[17]),
		.o_result(result14[2]), .o_cout(cout14[2]));
pu pu14_3 (.i_a(result13[2]), .i_b(~i_divisor[3]), .i_cin(cout14[2]), .i_carry_output(quotient[17]),
		.o_result(result14[3]), .o_cout(cout14[3]));
pu pu14_4 (.i_a(result13[3]), .i_b(~i_divisor[4]), .i_cin(cout14[3]), .i_carry_output(quotient[17]),
		.o_result(result14[4]), .o_cout(cout14[4]));
pu pu14_5 (.i_a(result13[4]), .i_b(~i_divisor[5]), .i_cin(cout14[4]), .i_carry_output(quotient[17]),
		.o_result(result14[5]), .o_cout(cout14[5]));
pu pu14_6 (.i_a(result13[5]), .i_b(~i_divisor[6]), .i_cin(cout14[5]), .i_carry_output(quotient[17]),
		.o_result(result14[6]), .o_cout(cout14[6]));
pu pu14_7 (.i_a(result13[6]), .i_b(~i_divisor[7]), .i_cin(cout14[6]), .i_carry_output(quotient[17]),
		.o_result(result14[7]), .o_cout(cout14[7]));
pu pu14_8 (.i_a(result13[7]), .i_b(~i_divisor[8]), .i_cin(cout14[7]), .i_carry_output(quotient[17]),
		.o_result(result14[8]), .o_cout(cout14[8]));
pu pu14_9 (.i_a(result13[8]), .i_b(~i_divisor[9]), .i_cin(cout14[8]), .i_carry_output(quotient[17]),
		.o_result(result14[9]), .o_cout(cout14[9]));
pu pu14_10 (.i_a(result13[9]), .i_b(~i_divisor[10]), .i_cin(cout14[9]), .i_carry_output(quotient[17]),
		.o_result(result14[10]), .o_cout(cout14[10]));
pu pu14_11 (.i_a(result13[10]), .i_b(~i_divisor[11]), .i_cin(cout14[10]), .i_carry_output(quotient[17]),
		.o_result(result14[11]), .o_cout(cout14[11]));
pu pu14_12 (.i_a(result13[11]), .i_b(~i_divisor[12]), .i_cin(cout14[11]), .i_carry_output(quotient[17]),
		.o_result(result14[12]), .o_cout(cout14[12]));
pu pu14_13 (.i_a(result13[12]), .i_b(~i_divisor[13]), .i_cin(cout14[12]), .i_carry_output(quotient[17]),
		.o_result(result14[13]), .o_cout(cout14[13]));
pu pu14_14 (.i_a(result13[13]), .i_b(~i_divisor[14]), .i_cin(cout14[13]), .i_carry_output(quotient[17]),
		.o_result(result14[14]), .o_cout(cout14[14]));
pu pu14_15 (.i_a(result13[14]), .i_b(~i_divisor[15]), .i_cin(cout14[14]), .i_carry_output(quotient[17]),
		.o_result(result14[15]), .o_cout(cout14[15]));
pu pu14_16 (.i_a(result13[15]), .i_b(~i_divisor[16]), .i_cin(cout14[15]), .i_carry_output(quotient[17]),
		.o_result(result14[16]), .o_cout(cout14[16]));
pu pu14_17 (.i_a(result13[16]), .i_b(~i_divisor[17]), .i_cin(cout14[16]), .i_carry_output(quotient[17]),
		.o_result(result14[17]), .o_cout(cout14[17]));
pu pu14_18 (.i_a(result13[17]), .i_b(~i_divisor[18]), .i_cin(cout14[17]), .i_carry_output(quotient[17]),
		.o_result(result14[18]), .o_cout(cout14[18]));
pu pu14_19 (.i_a(result13[18]), .i_b(~i_divisor[19]), .i_cin(cout14[18]), .i_carry_output(quotient[17]),
		.o_result(result14[19]), .o_cout(cout14[19]));
pu pu14_20 (.i_a(result13[19]), .i_b(~i_divisor[20]), .i_cin(cout14[19]), .i_carry_output(quotient[17]),
		.o_result(result14[20]), .o_cout(cout14[20]));
pu pu14_21 (.i_a(result13[20]), .i_b(~i_divisor[21]), .i_cin(cout14[20]), .i_carry_output(quotient[17]),
		.o_result(result14[21]), .o_cout(cout14[21]));
pu pu14_22 (.i_a(result13[21]), .i_b(~i_divisor[22]), .i_cin(cout14[21]), .i_carry_output(quotient[17]),
		.o_result(result14[22]), .o_cout(cout14[22]));
pu pu14_23 (.i_a(result13[22]), .i_b(~i_divisor[23]), .i_cin(cout14[22]), .i_carry_output(quotient[17]),
		.o_result(result14[23]), .o_cout(cout14[23]));
pu pu14_24 (.i_a(result13[23]), .i_b(~i_divisor[24]), .i_cin(cout14[23]), .i_carry_output(quotient[17]),
		.o_result(result14[24]), .o_cout(cout14[24]));
pu pu14_25 (.i_a(result13[24]), .i_b(~i_divisor[25]), .i_cin(cout14[24]), .i_carry_output(quotient[17]),
		.o_result(result14[25]), .o_cout(cout14[25]));
pu pu14_26 (.i_a(result13[25]), .i_b(~i_divisor[26]), .i_cin(cout14[25]), .i_carry_output(quotient[17]),
		.o_result(result14[26]), .o_cout(cout14[26]));
pu pu14_27 (.i_a(result13[26]), .i_b(~i_divisor[27]), .i_cin(cout14[26]), .i_carry_output(quotient[17]),
		.o_result(result14[27]), .o_cout(cout14[27]));
pu pu14_28 (.i_a(result13[27]), .i_b(~i_divisor[28]), .i_cin(cout14[27]), .i_carry_output(quotient[17]),
		.o_result(result14[28]), .o_cout(cout14[28]));
pu pu14_29 (.i_a(result13[28]), .i_b(~i_divisor[29]), .i_cin(cout14[28]), .i_carry_output(quotient[17]),
		.o_result(result14[29]), .o_cout(cout14[29]));
pu pu14_30 (.i_a(result13[29]), .i_b(~i_divisor[30]), .i_cin(cout14[29]), .i_carry_output(quotient[17]),
		.o_result(result14[30]), .o_cout(cout14[30]));
pu pu14_31 (.i_a(result13[30]), .i_b(~i_divisor[31]), .i_cin(cout14[30]), .i_carry_output(quotient[17]),
		.o_cout(quotient[17]));

// Row 15
pu pu15_0 (.i_a(i_dividend[16]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[16]),
         .o_result(result15[0]), .o_cout(cout15[0]));
pu pu15_1 (.i_a(result14[0]), .i_b(~i_divisor[1]), .i_cin(cout15[0]), .i_carry_output(quotient[16]),
		.o_result(result15[1]), .o_cout(cout15[1]));
pu pu15_2 (.i_a(result14[1]), .i_b(~i_divisor[2]), .i_cin(cout15[1]), .i_carry_output(quotient[16]),
		.o_result(result15[2]), .o_cout(cout15[2]));
pu pu15_3 (.i_a(result14[2]), .i_b(~i_divisor[3]), .i_cin(cout15[2]), .i_carry_output(quotient[16]),
		.o_result(result15[3]), .o_cout(cout15[3]));
pu pu15_4 (.i_a(result14[3]), .i_b(~i_divisor[4]), .i_cin(cout15[3]), .i_carry_output(quotient[16]),
		.o_result(result15[4]), .o_cout(cout15[4]));
pu pu15_5 (.i_a(result14[4]), .i_b(~i_divisor[5]), .i_cin(cout15[4]), .i_carry_output(quotient[16]),
		.o_result(result15[5]), .o_cout(cout15[5]));
pu pu15_6 (.i_a(result14[5]), .i_b(~i_divisor[6]), .i_cin(cout15[5]), .i_carry_output(quotient[16]),
		.o_result(result15[6]), .o_cout(cout15[6]));
pu pu15_7 (.i_a(result14[6]), .i_b(~i_divisor[7]), .i_cin(cout15[6]), .i_carry_output(quotient[16]),
		.o_result(result15[7]), .o_cout(cout15[7]));
pu pu15_8 (.i_a(result14[7]), .i_b(~i_divisor[8]), .i_cin(cout15[7]), .i_carry_output(quotient[16]),
		.o_result(result15[8]), .o_cout(cout15[8]));
pu pu15_9 (.i_a(result14[8]), .i_b(~i_divisor[9]), .i_cin(cout15[8]), .i_carry_output(quotient[16]),
		.o_result(result15[9]), .o_cout(cout15[9]));
pu pu15_10 (.i_a(result14[9]), .i_b(~i_divisor[10]), .i_cin(cout15[9]), .i_carry_output(quotient[16]),
		.o_result(result15[10]), .o_cout(cout15[10]));
pu pu15_11 (.i_a(result14[10]), .i_b(~i_divisor[11]), .i_cin(cout15[10]), .i_carry_output(quotient[16]),
		.o_result(result15[11]), .o_cout(cout15[11]));
pu pu15_12 (.i_a(result14[11]), .i_b(~i_divisor[12]), .i_cin(cout15[11]), .i_carry_output(quotient[16]),
		.o_result(result15[12]), .o_cout(cout15[12]));
pu pu15_13 (.i_a(result14[12]), .i_b(~i_divisor[13]), .i_cin(cout15[12]), .i_carry_output(quotient[16]),
		.o_result(result15[13]), .o_cout(cout15[13]));
pu pu15_14 (.i_a(result14[13]), .i_b(~i_divisor[14]), .i_cin(cout15[13]), .i_carry_output(quotient[16]),
		.o_result(result15[14]), .o_cout(cout15[14]));
pu pu15_15 (.i_a(result14[14]), .i_b(~i_divisor[15]), .i_cin(cout15[14]), .i_carry_output(quotient[16]),
		.o_result(result15[15]), .o_cout(cout15[15]));
pu pu15_16 (.i_a(result14[15]), .i_b(~i_divisor[16]), .i_cin(cout15[15]), .i_carry_output(quotient[16]),
		.o_result(result15[16]), .o_cout(cout15[16]));
pu pu15_17 (.i_a(result14[16]), .i_b(~i_divisor[17]), .i_cin(cout15[16]), .i_carry_output(quotient[16]),
		.o_result(result15[17]), .o_cout(cout15[17]));
pu pu15_18 (.i_a(result14[17]), .i_b(~i_divisor[18]), .i_cin(cout15[17]), .i_carry_output(quotient[16]),
		.o_result(result15[18]), .o_cout(cout15[18]));
pu pu15_19 (.i_a(result14[18]), .i_b(~i_divisor[19]), .i_cin(cout15[18]), .i_carry_output(quotient[16]),
		.o_result(result15[19]), .o_cout(cout15[19]));
pu pu15_20 (.i_a(result14[19]), .i_b(~i_divisor[20]), .i_cin(cout15[19]), .i_carry_output(quotient[16]),
		.o_result(result15[20]), .o_cout(cout15[20]));
pu pu15_21 (.i_a(result14[20]), .i_b(~i_divisor[21]), .i_cin(cout15[20]), .i_carry_output(quotient[16]),
		.o_result(result15[21]), .o_cout(cout15[21]));
pu pu15_22 (.i_a(result14[21]), .i_b(~i_divisor[22]), .i_cin(cout15[21]), .i_carry_output(quotient[16]),
		.o_result(result15[22]), .o_cout(cout15[22]));
pu pu15_23 (.i_a(result14[22]), .i_b(~i_divisor[23]), .i_cin(cout15[22]), .i_carry_output(quotient[16]),
		.o_result(result15[23]), .o_cout(cout15[23]));
pu pu15_24 (.i_a(result14[23]), .i_b(~i_divisor[24]), .i_cin(cout15[23]), .i_carry_output(quotient[16]),
		.o_result(result15[24]), .o_cout(cout15[24]));
pu pu15_25 (.i_a(result14[24]), .i_b(~i_divisor[25]), .i_cin(cout15[24]), .i_carry_output(quotient[16]),
		.o_result(result15[25]), .o_cout(cout15[25]));
pu pu15_26 (.i_a(result14[25]), .i_b(~i_divisor[26]), .i_cin(cout15[25]), .i_carry_output(quotient[16]),
		.o_result(result15[26]), .o_cout(cout15[26]));
pu pu15_27 (.i_a(result14[26]), .i_b(~i_divisor[27]), .i_cin(cout15[26]), .i_carry_output(quotient[16]),
		.o_result(result15[27]), .o_cout(cout15[27]));
pu pu15_28 (.i_a(result14[27]), .i_b(~i_divisor[28]), .i_cin(cout15[27]), .i_carry_output(quotient[16]),
		.o_result(result15[28]), .o_cout(cout15[28]));
pu pu15_29 (.i_a(result14[28]), .i_b(~i_divisor[29]), .i_cin(cout15[28]), .i_carry_output(quotient[16]),
		.o_result(result15[29]), .o_cout(cout15[29]));
pu pu15_30 (.i_a(result14[29]), .i_b(~i_divisor[30]), .i_cin(cout15[29]), .i_carry_output(quotient[16]),
		.o_result(result15[30]), .o_cout(cout15[30]));
pu pu15_31 (.i_a(result14[30]), .i_b(~i_divisor[31]), .i_cin(cout15[30]), .i_carry_output(quotient[16]),
		.o_cout(quotient[16]));

// Row 16
pu pu16_0 (.i_a(i_dividend[15]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[15]),
         .o_result(result16[0]), .o_cout(cout16[0]));
pu pu16_1 (.i_a(result15[0]), .i_b(~i_divisor[1]), .i_cin(cout16[0]), .i_carry_output(quotient[15]),
		.o_result(result16[1]), .o_cout(cout16[1]));
pu pu16_2 (.i_a(result15[1]), .i_b(~i_divisor[2]), .i_cin(cout16[1]), .i_carry_output(quotient[15]),
		.o_result(result16[2]), .o_cout(cout16[2]));
pu pu16_3 (.i_a(result15[2]), .i_b(~i_divisor[3]), .i_cin(cout16[2]), .i_carry_output(quotient[15]),
		.o_result(result16[3]), .o_cout(cout16[3]));
pu pu16_4 (.i_a(result15[3]), .i_b(~i_divisor[4]), .i_cin(cout16[3]), .i_carry_output(quotient[15]),
		.o_result(result16[4]), .o_cout(cout16[4]));
pu pu16_5 (.i_a(result15[4]), .i_b(~i_divisor[5]), .i_cin(cout16[4]), .i_carry_output(quotient[15]),
		.o_result(result16[5]), .o_cout(cout16[5]));
pu pu16_6 (.i_a(result15[5]), .i_b(~i_divisor[6]), .i_cin(cout16[5]), .i_carry_output(quotient[15]),
		.o_result(result16[6]), .o_cout(cout16[6]));
pu pu16_7 (.i_a(result15[6]), .i_b(~i_divisor[7]), .i_cin(cout16[6]), .i_carry_output(quotient[15]),
		.o_result(result16[7]), .o_cout(cout16[7]));
pu pu16_8 (.i_a(result15[7]), .i_b(~i_divisor[8]), .i_cin(cout16[7]), .i_carry_output(quotient[15]),
		.o_result(result16[8]), .o_cout(cout16[8]));
pu pu16_9 (.i_a(result15[8]), .i_b(~i_divisor[9]), .i_cin(cout16[8]), .i_carry_output(quotient[15]),
		.o_result(result16[9]), .o_cout(cout16[9]));
pu pu16_10 (.i_a(result15[9]), .i_b(~i_divisor[10]), .i_cin(cout16[9]), .i_carry_output(quotient[15]),
		.o_result(result16[10]), .o_cout(cout16[10]));
pu pu16_11 (.i_a(result15[10]), .i_b(~i_divisor[11]), .i_cin(cout16[10]), .i_carry_output(quotient[15]),
		.o_result(result16[11]), .o_cout(cout16[11]));
pu pu16_12 (.i_a(result15[11]), .i_b(~i_divisor[12]), .i_cin(cout16[11]), .i_carry_output(quotient[15]),
		.o_result(result16[12]), .o_cout(cout16[12]));
pu pu16_13 (.i_a(result15[12]), .i_b(~i_divisor[13]), .i_cin(cout16[12]), .i_carry_output(quotient[15]),
		.o_result(result16[13]), .o_cout(cout16[13]));
pu pu16_14 (.i_a(result15[13]), .i_b(~i_divisor[14]), .i_cin(cout16[13]), .i_carry_output(quotient[15]),
		.o_result(result16[14]), .o_cout(cout16[14]));
pu pu16_15 (.i_a(result15[14]), .i_b(~i_divisor[15]), .i_cin(cout16[14]), .i_carry_output(quotient[15]),
		.o_result(result16[15]), .o_cout(cout16[15]));
pu pu16_16 (.i_a(result15[15]), .i_b(~i_divisor[16]), .i_cin(cout16[15]), .i_carry_output(quotient[15]),
		.o_result(result16[16]), .o_cout(cout16[16]));
pu pu16_17 (.i_a(result15[16]), .i_b(~i_divisor[17]), .i_cin(cout16[16]), .i_carry_output(quotient[15]),
		.o_result(result16[17]), .o_cout(cout16[17]));
pu pu16_18 (.i_a(result15[17]), .i_b(~i_divisor[18]), .i_cin(cout16[17]), .i_carry_output(quotient[15]),
		.o_result(result16[18]), .o_cout(cout16[18]));
pu pu16_19 (.i_a(result15[18]), .i_b(~i_divisor[19]), .i_cin(cout16[18]), .i_carry_output(quotient[15]),
		.o_result(result16[19]), .o_cout(cout16[19]));
pu pu16_20 (.i_a(result15[19]), .i_b(~i_divisor[20]), .i_cin(cout16[19]), .i_carry_output(quotient[15]),
		.o_result(result16[20]), .o_cout(cout16[20]));
pu pu16_21 (.i_a(result15[20]), .i_b(~i_divisor[21]), .i_cin(cout16[20]), .i_carry_output(quotient[15]),
		.o_result(result16[21]), .o_cout(cout16[21]));
pu pu16_22 (.i_a(result15[21]), .i_b(~i_divisor[22]), .i_cin(cout16[21]), .i_carry_output(quotient[15]),
		.o_result(result16[22]), .o_cout(cout16[22]));
pu pu16_23 (.i_a(result15[22]), .i_b(~i_divisor[23]), .i_cin(cout16[22]), .i_carry_output(quotient[15]),
		.o_result(result16[23]), .o_cout(cout16[23]));
pu pu16_24 (.i_a(result15[23]), .i_b(~i_divisor[24]), .i_cin(cout16[23]), .i_carry_output(quotient[15]),
		.o_result(result16[24]), .o_cout(cout16[24]));
pu pu16_25 (.i_a(result15[24]), .i_b(~i_divisor[25]), .i_cin(cout16[24]), .i_carry_output(quotient[15]),
		.o_result(result16[25]), .o_cout(cout16[25]));
pu pu16_26 (.i_a(result15[25]), .i_b(~i_divisor[26]), .i_cin(cout16[25]), .i_carry_output(quotient[15]),
		.o_result(result16[26]), .o_cout(cout16[26]));
pu pu16_27 (.i_a(result15[26]), .i_b(~i_divisor[27]), .i_cin(cout16[26]), .i_carry_output(quotient[15]),
		.o_result(result16[27]), .o_cout(cout16[27]));
pu pu16_28 (.i_a(result15[27]), .i_b(~i_divisor[28]), .i_cin(cout16[27]), .i_carry_output(quotient[15]),
		.o_result(result16[28]), .o_cout(cout16[28]));
pu pu16_29 (.i_a(result15[28]), .i_b(~i_divisor[29]), .i_cin(cout16[28]), .i_carry_output(quotient[15]),
		.o_result(result16[29]), .o_cout(cout16[29]));
pu pu16_30 (.i_a(result15[29]), .i_b(~i_divisor[30]), .i_cin(cout16[29]), .i_carry_output(quotient[15]),
		.o_result(result16[30]), .o_cout(cout16[30]));
pu pu16_31 (.i_a(result15[30]), .i_b(~i_divisor[31]), .i_cin(cout16[30]), .i_carry_output(quotient[15]),
		.o_cout(quotient[15]));

// Row 17
pu pu17_0 (.i_a(i_dividend[14]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[14]),
         .o_result(result17[0]), .o_cout(cout17[0]));
pu pu17_1 (.i_a(result16[0]), .i_b(~i_divisor[1]), .i_cin(cout17[0]), .i_carry_output(quotient[14]),
		.o_result(result17[1]), .o_cout(cout17[1]));
pu pu17_2 (.i_a(result16[1]), .i_b(~i_divisor[2]), .i_cin(cout17[1]), .i_carry_output(quotient[14]),
		.o_result(result17[2]), .o_cout(cout17[2]));
pu pu17_3 (.i_a(result16[2]), .i_b(~i_divisor[3]), .i_cin(cout17[2]), .i_carry_output(quotient[14]),
		.o_result(result17[3]), .o_cout(cout17[3]));
pu pu17_4 (.i_a(result16[3]), .i_b(~i_divisor[4]), .i_cin(cout17[3]), .i_carry_output(quotient[14]),
		.o_result(result17[4]), .o_cout(cout17[4]));
pu pu17_5 (.i_a(result16[4]), .i_b(~i_divisor[5]), .i_cin(cout17[4]), .i_carry_output(quotient[14]),
		.o_result(result17[5]), .o_cout(cout17[5]));
pu pu17_6 (.i_a(result16[5]), .i_b(~i_divisor[6]), .i_cin(cout17[5]), .i_carry_output(quotient[14]),
		.o_result(result17[6]), .o_cout(cout17[6]));
pu pu17_7 (.i_a(result16[6]), .i_b(~i_divisor[7]), .i_cin(cout17[6]), .i_carry_output(quotient[14]),
		.o_result(result17[7]), .o_cout(cout17[7]));
pu pu17_8 (.i_a(result16[7]), .i_b(~i_divisor[8]), .i_cin(cout17[7]), .i_carry_output(quotient[14]),
		.o_result(result17[8]), .o_cout(cout17[8]));
pu pu17_9 (.i_a(result16[8]), .i_b(~i_divisor[9]), .i_cin(cout17[8]), .i_carry_output(quotient[14]),
		.o_result(result17[9]), .o_cout(cout17[9]));
pu pu17_10 (.i_a(result16[9]), .i_b(~i_divisor[10]), .i_cin(cout17[9]), .i_carry_output(quotient[14]),
		.o_result(result17[10]), .o_cout(cout17[10]));
pu pu17_11 (.i_a(result16[10]), .i_b(~i_divisor[11]), .i_cin(cout17[10]), .i_carry_output(quotient[14]),
		.o_result(result17[11]), .o_cout(cout17[11]));
pu pu17_12 (.i_a(result16[11]), .i_b(~i_divisor[12]), .i_cin(cout17[11]), .i_carry_output(quotient[14]),
		.o_result(result17[12]), .o_cout(cout17[12]));
pu pu17_13 (.i_a(result16[12]), .i_b(~i_divisor[13]), .i_cin(cout17[12]), .i_carry_output(quotient[14]),
		.o_result(result17[13]), .o_cout(cout17[13]));
pu pu17_14 (.i_a(result16[13]), .i_b(~i_divisor[14]), .i_cin(cout17[13]), .i_carry_output(quotient[14]),
		.o_result(result17[14]), .o_cout(cout17[14]));
pu pu17_15 (.i_a(result16[14]), .i_b(~i_divisor[15]), .i_cin(cout17[14]), .i_carry_output(quotient[14]),
		.o_result(result17[15]), .o_cout(cout17[15]));
pu pu17_16 (.i_a(result16[15]), .i_b(~i_divisor[16]), .i_cin(cout17[15]), .i_carry_output(quotient[14]),
		.o_result(result17[16]), .o_cout(cout17[16]));
pu pu17_17 (.i_a(result16[16]), .i_b(~i_divisor[17]), .i_cin(cout17[16]), .i_carry_output(quotient[14]),
		.o_result(result17[17]), .o_cout(cout17[17]));
pu pu17_18 (.i_a(result16[17]), .i_b(~i_divisor[18]), .i_cin(cout17[17]), .i_carry_output(quotient[14]),
		.o_result(result17[18]), .o_cout(cout17[18]));
pu pu17_19 (.i_a(result16[18]), .i_b(~i_divisor[19]), .i_cin(cout17[18]), .i_carry_output(quotient[14]),
		.o_result(result17[19]), .o_cout(cout17[19]));
pu pu17_20 (.i_a(result16[19]), .i_b(~i_divisor[20]), .i_cin(cout17[19]), .i_carry_output(quotient[14]),
		.o_result(result17[20]), .o_cout(cout17[20]));
pu pu17_21 (.i_a(result16[20]), .i_b(~i_divisor[21]), .i_cin(cout17[20]), .i_carry_output(quotient[14]),
		.o_result(result17[21]), .o_cout(cout17[21]));
pu pu17_22 (.i_a(result16[21]), .i_b(~i_divisor[22]), .i_cin(cout17[21]), .i_carry_output(quotient[14]),
		.o_result(result17[22]), .o_cout(cout17[22]));
pu pu17_23 (.i_a(result16[22]), .i_b(~i_divisor[23]), .i_cin(cout17[22]), .i_carry_output(quotient[14]),
		.o_result(result17[23]), .o_cout(cout17[23]));
pu pu17_24 (.i_a(result16[23]), .i_b(~i_divisor[24]), .i_cin(cout17[23]), .i_carry_output(quotient[14]),
		.o_result(result17[24]), .o_cout(cout17[24]));
pu pu17_25 (.i_a(result16[24]), .i_b(~i_divisor[25]), .i_cin(cout17[24]), .i_carry_output(quotient[14]),
		.o_result(result17[25]), .o_cout(cout17[25]));
pu pu17_26 (.i_a(result16[25]), .i_b(~i_divisor[26]), .i_cin(cout17[25]), .i_carry_output(quotient[14]),
		.o_result(result17[26]), .o_cout(cout17[26]));
pu pu17_27 (.i_a(result16[26]), .i_b(~i_divisor[27]), .i_cin(cout17[26]), .i_carry_output(quotient[14]),
		.o_result(result17[27]), .o_cout(cout17[27]));
pu pu17_28 (.i_a(result16[27]), .i_b(~i_divisor[28]), .i_cin(cout17[27]), .i_carry_output(quotient[14]),
		.o_result(result17[28]), .o_cout(cout17[28]));
pu pu17_29 (.i_a(result16[28]), .i_b(~i_divisor[29]), .i_cin(cout17[28]), .i_carry_output(quotient[14]),
		.o_result(result17[29]), .o_cout(cout17[29]));
pu pu17_30 (.i_a(result16[29]), .i_b(~i_divisor[30]), .i_cin(cout17[29]), .i_carry_output(quotient[14]),
		.o_result(result17[30]), .o_cout(cout17[30]));
pu pu17_31 (.i_a(result16[30]), .i_b(~i_divisor[31]), .i_cin(cout17[30]), .i_carry_output(quotient[14]),
		.o_cout(quotient[14]));

// Row 18
pu pu18_0 (.i_a(i_dividend[13]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[13]),
         .o_result(result18[0]), .o_cout(cout18[0]));
pu pu18_1 (.i_a(result17[0]), .i_b(~i_divisor[1]), .i_cin(cout18[0]), .i_carry_output(quotient[13]),
		.o_result(result18[1]), .o_cout(cout18[1]));
pu pu18_2 (.i_a(result17[1]), .i_b(~i_divisor[2]), .i_cin(cout18[1]), .i_carry_output(quotient[13]),
		.o_result(result18[2]), .o_cout(cout18[2]));
pu pu18_3 (.i_a(result17[2]), .i_b(~i_divisor[3]), .i_cin(cout18[2]), .i_carry_output(quotient[13]),
		.o_result(result18[3]), .o_cout(cout18[3]));
pu pu18_4 (.i_a(result17[3]), .i_b(~i_divisor[4]), .i_cin(cout18[3]), .i_carry_output(quotient[13]),
		.o_result(result18[4]), .o_cout(cout18[4]));
pu pu18_5 (.i_a(result17[4]), .i_b(~i_divisor[5]), .i_cin(cout18[4]), .i_carry_output(quotient[13]),
		.o_result(result18[5]), .o_cout(cout18[5]));
pu pu18_6 (.i_a(result17[5]), .i_b(~i_divisor[6]), .i_cin(cout18[5]), .i_carry_output(quotient[13]),
		.o_result(result18[6]), .o_cout(cout18[6]));
pu pu18_7 (.i_a(result17[6]), .i_b(~i_divisor[7]), .i_cin(cout18[6]), .i_carry_output(quotient[13]),
		.o_result(result18[7]), .o_cout(cout18[7]));
pu pu18_8 (.i_a(result17[7]), .i_b(~i_divisor[8]), .i_cin(cout18[7]), .i_carry_output(quotient[13]),
		.o_result(result18[8]), .o_cout(cout18[8]));
pu pu18_9 (.i_a(result17[8]), .i_b(~i_divisor[9]), .i_cin(cout18[8]), .i_carry_output(quotient[13]),
		.o_result(result18[9]), .o_cout(cout18[9]));
pu pu18_10 (.i_a(result17[9]), .i_b(~i_divisor[10]), .i_cin(cout18[9]), .i_carry_output(quotient[13]),
		.o_result(result18[10]), .o_cout(cout18[10]));
pu pu18_11 (.i_a(result17[10]), .i_b(~i_divisor[11]), .i_cin(cout18[10]), .i_carry_output(quotient[13]),
		.o_result(result18[11]), .o_cout(cout18[11]));
pu pu18_12 (.i_a(result17[11]), .i_b(~i_divisor[12]), .i_cin(cout18[11]), .i_carry_output(quotient[13]),
		.o_result(result18[12]), .o_cout(cout18[12]));
pu pu18_13 (.i_a(result17[12]), .i_b(~i_divisor[13]), .i_cin(cout18[12]), .i_carry_output(quotient[13]),
		.o_result(result18[13]), .o_cout(cout18[13]));
pu pu18_14 (.i_a(result17[13]), .i_b(~i_divisor[14]), .i_cin(cout18[13]), .i_carry_output(quotient[13]),
		.o_result(result18[14]), .o_cout(cout18[14]));
pu pu18_15 (.i_a(result17[14]), .i_b(~i_divisor[15]), .i_cin(cout18[14]), .i_carry_output(quotient[13]),
		.o_result(result18[15]), .o_cout(cout18[15]));
pu pu18_16 (.i_a(result17[15]), .i_b(~i_divisor[16]), .i_cin(cout18[15]), .i_carry_output(quotient[13]),
		.o_result(result18[16]), .o_cout(cout18[16]));
pu pu18_17 (.i_a(result17[16]), .i_b(~i_divisor[17]), .i_cin(cout18[16]), .i_carry_output(quotient[13]),
		.o_result(result18[17]), .o_cout(cout18[17]));
pu pu18_18 (.i_a(result17[17]), .i_b(~i_divisor[18]), .i_cin(cout18[17]), .i_carry_output(quotient[13]),
		.o_result(result18[18]), .o_cout(cout18[18]));
pu pu18_19 (.i_a(result17[18]), .i_b(~i_divisor[19]), .i_cin(cout18[18]), .i_carry_output(quotient[13]),
		.o_result(result18[19]), .o_cout(cout18[19]));
pu pu18_20 (.i_a(result17[19]), .i_b(~i_divisor[20]), .i_cin(cout18[19]), .i_carry_output(quotient[13]),
		.o_result(result18[20]), .o_cout(cout18[20]));
pu pu18_21 (.i_a(result17[20]), .i_b(~i_divisor[21]), .i_cin(cout18[20]), .i_carry_output(quotient[13]),
		.o_result(result18[21]), .o_cout(cout18[21]));
pu pu18_22 (.i_a(result17[21]), .i_b(~i_divisor[22]), .i_cin(cout18[21]), .i_carry_output(quotient[13]),
		.o_result(result18[22]), .o_cout(cout18[22]));
pu pu18_23 (.i_a(result17[22]), .i_b(~i_divisor[23]), .i_cin(cout18[22]), .i_carry_output(quotient[13]),
		.o_result(result18[23]), .o_cout(cout18[23]));
pu pu18_24 (.i_a(result17[23]), .i_b(~i_divisor[24]), .i_cin(cout18[23]), .i_carry_output(quotient[13]),
		.o_result(result18[24]), .o_cout(cout18[24]));
pu pu18_25 (.i_a(result17[24]), .i_b(~i_divisor[25]), .i_cin(cout18[24]), .i_carry_output(quotient[13]),
		.o_result(result18[25]), .o_cout(cout18[25]));
pu pu18_26 (.i_a(result17[25]), .i_b(~i_divisor[26]), .i_cin(cout18[25]), .i_carry_output(quotient[13]),
		.o_result(result18[26]), .o_cout(cout18[26]));
pu pu18_27 (.i_a(result17[26]), .i_b(~i_divisor[27]), .i_cin(cout18[26]), .i_carry_output(quotient[13]),
		.o_result(result18[27]), .o_cout(cout18[27]));
pu pu18_28 (.i_a(result17[27]), .i_b(~i_divisor[28]), .i_cin(cout18[27]), .i_carry_output(quotient[13]),
		.o_result(result18[28]), .o_cout(cout18[28]));
pu pu18_29 (.i_a(result17[28]), .i_b(~i_divisor[29]), .i_cin(cout18[28]), .i_carry_output(quotient[13]),
		.o_result(result18[29]), .o_cout(cout18[29]));
pu pu18_30 (.i_a(result17[29]), .i_b(~i_divisor[30]), .i_cin(cout18[29]), .i_carry_output(quotient[13]),
		.o_result(result18[30]), .o_cout(cout18[30]));
pu pu18_31 (.i_a(result17[30]), .i_b(~i_divisor[31]), .i_cin(cout18[30]), .i_carry_output(quotient[13]),
		.o_cout(quotient[13]));

// Row 19
pu pu19_0 (.i_a(i_dividend[12]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[12]),
         .o_result(result19[0]), .o_cout(cout19[0]));
pu pu19_1 (.i_a(result18[0]), .i_b(~i_divisor[1]), .i_cin(cout19[0]), .i_carry_output(quotient[12]),
		.o_result(result19[1]), .o_cout(cout19[1]));
pu pu19_2 (.i_a(result18[1]), .i_b(~i_divisor[2]), .i_cin(cout19[1]), .i_carry_output(quotient[12]),
		.o_result(result19[2]), .o_cout(cout19[2]));
pu pu19_3 (.i_a(result18[2]), .i_b(~i_divisor[3]), .i_cin(cout19[2]), .i_carry_output(quotient[12]),
		.o_result(result19[3]), .o_cout(cout19[3]));
pu pu19_4 (.i_a(result18[3]), .i_b(~i_divisor[4]), .i_cin(cout19[3]), .i_carry_output(quotient[12]),
		.o_result(result19[4]), .o_cout(cout19[4]));
pu pu19_5 (.i_a(result18[4]), .i_b(~i_divisor[5]), .i_cin(cout19[4]), .i_carry_output(quotient[12]),
		.o_result(result19[5]), .o_cout(cout19[5]));
pu pu19_6 (.i_a(result18[5]), .i_b(~i_divisor[6]), .i_cin(cout19[5]), .i_carry_output(quotient[12]),
		.o_result(result19[6]), .o_cout(cout19[6]));
pu pu19_7 (.i_a(result18[6]), .i_b(~i_divisor[7]), .i_cin(cout19[6]), .i_carry_output(quotient[12]),
		.o_result(result19[7]), .o_cout(cout19[7]));
pu pu19_8 (.i_a(result18[7]), .i_b(~i_divisor[8]), .i_cin(cout19[7]), .i_carry_output(quotient[12]),
		.o_result(result19[8]), .o_cout(cout19[8]));
pu pu19_9 (.i_a(result18[8]), .i_b(~i_divisor[9]), .i_cin(cout19[8]), .i_carry_output(quotient[12]),
		.o_result(result19[9]), .o_cout(cout19[9]));
pu pu19_10 (.i_a(result18[9]), .i_b(~i_divisor[10]), .i_cin(cout19[9]), .i_carry_output(quotient[12]),
		.o_result(result19[10]), .o_cout(cout19[10]));
pu pu19_11 (.i_a(result18[10]), .i_b(~i_divisor[11]), .i_cin(cout19[10]), .i_carry_output(quotient[12]),
		.o_result(result19[11]), .o_cout(cout19[11]));
pu pu19_12 (.i_a(result18[11]), .i_b(~i_divisor[12]), .i_cin(cout19[11]), .i_carry_output(quotient[12]),
		.o_result(result19[12]), .o_cout(cout19[12]));
pu pu19_13 (.i_a(result18[12]), .i_b(~i_divisor[13]), .i_cin(cout19[12]), .i_carry_output(quotient[12]),
		.o_result(result19[13]), .o_cout(cout19[13]));
pu pu19_14 (.i_a(result18[13]), .i_b(~i_divisor[14]), .i_cin(cout19[13]), .i_carry_output(quotient[12]),
		.o_result(result19[14]), .o_cout(cout19[14]));
pu pu19_15 (.i_a(result18[14]), .i_b(~i_divisor[15]), .i_cin(cout19[14]), .i_carry_output(quotient[12]),
		.o_result(result19[15]), .o_cout(cout19[15]));
pu pu19_16 (.i_a(result18[15]), .i_b(~i_divisor[16]), .i_cin(cout19[15]), .i_carry_output(quotient[12]),
		.o_result(result19[16]), .o_cout(cout19[16]));
pu pu19_17 (.i_a(result18[16]), .i_b(~i_divisor[17]), .i_cin(cout19[16]), .i_carry_output(quotient[12]),
		.o_result(result19[17]), .o_cout(cout19[17]));
pu pu19_18 (.i_a(result18[17]), .i_b(~i_divisor[18]), .i_cin(cout19[17]), .i_carry_output(quotient[12]),
		.o_result(result19[18]), .o_cout(cout19[18]));
pu pu19_19 (.i_a(result18[18]), .i_b(~i_divisor[19]), .i_cin(cout19[18]), .i_carry_output(quotient[12]),
		.o_result(result19[19]), .o_cout(cout19[19]));
pu pu19_20 (.i_a(result18[19]), .i_b(~i_divisor[20]), .i_cin(cout19[19]), .i_carry_output(quotient[12]),
		.o_result(result19[20]), .o_cout(cout19[20]));
pu pu19_21 (.i_a(result18[20]), .i_b(~i_divisor[21]), .i_cin(cout19[20]), .i_carry_output(quotient[12]),
		.o_result(result19[21]), .o_cout(cout19[21]));
pu pu19_22 (.i_a(result18[21]), .i_b(~i_divisor[22]), .i_cin(cout19[21]), .i_carry_output(quotient[12]),
		.o_result(result19[22]), .o_cout(cout19[22]));
pu pu19_23 (.i_a(result18[22]), .i_b(~i_divisor[23]), .i_cin(cout19[22]), .i_carry_output(quotient[12]),
		.o_result(result19[23]), .o_cout(cout19[23]));
pu pu19_24 (.i_a(result18[23]), .i_b(~i_divisor[24]), .i_cin(cout19[23]), .i_carry_output(quotient[12]),
		.o_result(result19[24]), .o_cout(cout19[24]));
pu pu19_25 (.i_a(result18[24]), .i_b(~i_divisor[25]), .i_cin(cout19[24]), .i_carry_output(quotient[12]),
		.o_result(result19[25]), .o_cout(cout19[25]));
pu pu19_26 (.i_a(result18[25]), .i_b(~i_divisor[26]), .i_cin(cout19[25]), .i_carry_output(quotient[12]),
		.o_result(result19[26]), .o_cout(cout19[26]));
pu pu19_27 (.i_a(result18[26]), .i_b(~i_divisor[27]), .i_cin(cout19[26]), .i_carry_output(quotient[12]),
		.o_result(result19[27]), .o_cout(cout19[27]));
pu pu19_28 (.i_a(result18[27]), .i_b(~i_divisor[28]), .i_cin(cout19[27]), .i_carry_output(quotient[12]),
		.o_result(result19[28]), .o_cout(cout19[28]));
pu pu19_29 (.i_a(result18[28]), .i_b(~i_divisor[29]), .i_cin(cout19[28]), .i_carry_output(quotient[12]),
		.o_result(result19[29]), .o_cout(cout19[29]));
pu pu19_30 (.i_a(result18[29]), .i_b(~i_divisor[30]), .i_cin(cout19[29]), .i_carry_output(quotient[12]),
		.o_result(result19[30]), .o_cout(cout19[30]));
pu pu19_31 (.i_a(result18[30]), .i_b(~i_divisor[31]), .i_cin(cout19[30]), .i_carry_output(quotient[12]),
		.o_cout(quotient[12]));

// Row 20
pu pu20_0 (.i_a(i_dividend[11]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[11]),
         .o_result(result20[0]), .o_cout(cout20[0]));
pu pu20_1 (.i_a(result19[0]), .i_b(~i_divisor[1]), .i_cin(cout20[0]), .i_carry_output(quotient[11]),
		.o_result(result20[1]), .o_cout(cout20[1]));
pu pu20_2 (.i_a(result19[1]), .i_b(~i_divisor[2]), .i_cin(cout20[1]), .i_carry_output(quotient[11]),
		.o_result(result20[2]), .o_cout(cout20[2]));
pu pu20_3 (.i_a(result19[2]), .i_b(~i_divisor[3]), .i_cin(cout20[2]), .i_carry_output(quotient[11]),
		.o_result(result20[3]), .o_cout(cout20[3]));
pu pu20_4 (.i_a(result19[3]), .i_b(~i_divisor[4]), .i_cin(cout20[3]), .i_carry_output(quotient[11]),
		.o_result(result20[4]), .o_cout(cout20[4]));
pu pu20_5 (.i_a(result19[4]), .i_b(~i_divisor[5]), .i_cin(cout20[4]), .i_carry_output(quotient[11]),
		.o_result(result20[5]), .o_cout(cout20[5]));
pu pu20_6 (.i_a(result19[5]), .i_b(~i_divisor[6]), .i_cin(cout20[5]), .i_carry_output(quotient[11]),
		.o_result(result20[6]), .o_cout(cout20[6]));
pu pu20_7 (.i_a(result19[6]), .i_b(~i_divisor[7]), .i_cin(cout20[6]), .i_carry_output(quotient[11]),
		.o_result(result20[7]), .o_cout(cout20[7]));
pu pu20_8 (.i_a(result19[7]), .i_b(~i_divisor[8]), .i_cin(cout20[7]), .i_carry_output(quotient[11]),
		.o_result(result20[8]), .o_cout(cout20[8]));
pu pu20_9 (.i_a(result19[8]), .i_b(~i_divisor[9]), .i_cin(cout20[8]), .i_carry_output(quotient[11]),
		.o_result(result20[9]), .o_cout(cout20[9]));
pu pu20_10 (.i_a(result19[9]), .i_b(~i_divisor[10]), .i_cin(cout20[9]), .i_carry_output(quotient[11]),
		.o_result(result20[10]), .o_cout(cout20[10]));
pu pu20_11 (.i_a(result19[10]), .i_b(~i_divisor[11]), .i_cin(cout20[10]), .i_carry_output(quotient[11]),
		.o_result(result20[11]), .o_cout(cout20[11]));
pu pu20_12 (.i_a(result19[11]), .i_b(~i_divisor[12]), .i_cin(cout20[11]), .i_carry_output(quotient[11]),
		.o_result(result20[12]), .o_cout(cout20[12]));
pu pu20_13 (.i_a(result19[12]), .i_b(~i_divisor[13]), .i_cin(cout20[12]), .i_carry_output(quotient[11]),
		.o_result(result20[13]), .o_cout(cout20[13]));
pu pu20_14 (.i_a(result19[13]), .i_b(~i_divisor[14]), .i_cin(cout20[13]), .i_carry_output(quotient[11]),
		.o_result(result20[14]), .o_cout(cout20[14]));
pu pu20_15 (.i_a(result19[14]), .i_b(~i_divisor[15]), .i_cin(cout20[14]), .i_carry_output(quotient[11]),
		.o_result(result20[15]), .o_cout(cout20[15]));
pu pu20_16 (.i_a(result19[15]), .i_b(~i_divisor[16]), .i_cin(cout20[15]), .i_carry_output(quotient[11]),
		.o_result(result20[16]), .o_cout(cout20[16]));
pu pu20_17 (.i_a(result19[16]), .i_b(~i_divisor[17]), .i_cin(cout20[16]), .i_carry_output(quotient[11]),
		.o_result(result20[17]), .o_cout(cout20[17]));
pu pu20_18 (.i_a(result19[17]), .i_b(~i_divisor[18]), .i_cin(cout20[17]), .i_carry_output(quotient[11]),
		.o_result(result20[18]), .o_cout(cout20[18]));
pu pu20_19 (.i_a(result19[18]), .i_b(~i_divisor[19]), .i_cin(cout20[18]), .i_carry_output(quotient[11]),
		.o_result(result20[19]), .o_cout(cout20[19]));
pu pu20_20 (.i_a(result19[19]), .i_b(~i_divisor[20]), .i_cin(cout20[19]), .i_carry_output(quotient[11]),
		.o_result(result20[20]), .o_cout(cout20[20]));
pu pu20_21 (.i_a(result19[20]), .i_b(~i_divisor[21]), .i_cin(cout20[20]), .i_carry_output(quotient[11]),
		.o_result(result20[21]), .o_cout(cout20[21]));
pu pu20_22 (.i_a(result19[21]), .i_b(~i_divisor[22]), .i_cin(cout20[21]), .i_carry_output(quotient[11]),
		.o_result(result20[22]), .o_cout(cout20[22]));
pu pu20_23 (.i_a(result19[22]), .i_b(~i_divisor[23]), .i_cin(cout20[22]), .i_carry_output(quotient[11]),
		.o_result(result20[23]), .o_cout(cout20[23]));
pu pu20_24 (.i_a(result19[23]), .i_b(~i_divisor[24]), .i_cin(cout20[23]), .i_carry_output(quotient[11]),
		.o_result(result20[24]), .o_cout(cout20[24]));
pu pu20_25 (.i_a(result19[24]), .i_b(~i_divisor[25]), .i_cin(cout20[24]), .i_carry_output(quotient[11]),
		.o_result(result20[25]), .o_cout(cout20[25]));
pu pu20_26 (.i_a(result19[25]), .i_b(~i_divisor[26]), .i_cin(cout20[25]), .i_carry_output(quotient[11]),
		.o_result(result20[26]), .o_cout(cout20[26]));
pu pu20_27 (.i_a(result19[26]), .i_b(~i_divisor[27]), .i_cin(cout20[26]), .i_carry_output(quotient[11]),
		.o_result(result20[27]), .o_cout(cout20[27]));
pu pu20_28 (.i_a(result19[27]), .i_b(~i_divisor[28]), .i_cin(cout20[27]), .i_carry_output(quotient[11]),
		.o_result(result20[28]), .o_cout(cout20[28]));
pu pu20_29 (.i_a(result19[28]), .i_b(~i_divisor[29]), .i_cin(cout20[28]), .i_carry_output(quotient[11]),
		.o_result(result20[29]), .o_cout(cout20[29]));
pu pu20_30 (.i_a(result19[29]), .i_b(~i_divisor[30]), .i_cin(cout20[29]), .i_carry_output(quotient[11]),
		.o_result(result20[30]), .o_cout(cout20[30]));
pu pu20_31 (.i_a(result19[30]), .i_b(~i_divisor[31]), .i_cin(cout20[30]), .i_carry_output(quotient[11]),
		.o_cout(quotient[11]));
		
// Row 21
pu pu21_0 (.i_a(i_dividend[10]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[10]),
         .o_result(result21[0]), .o_cout(cout21[0]));
pu pu21_1 (.i_a(result20[0]), .i_b(~i_divisor[1]), .i_cin(cout21[0]), .i_carry_output(quotient[10]),
		.o_result(result21[1]), .o_cout(cout21[1]));
pu pu21_2 (.i_a(result20[1]), .i_b(~i_divisor[2]), .i_cin(cout21[1]), .i_carry_output(quotient[10]),
		.o_result(result21[2]), .o_cout(cout21[2]));
pu pu21_3 (.i_a(result20[2]), .i_b(~i_divisor[3]), .i_cin(cout21[2]), .i_carry_output(quotient[10]),
		.o_result(result21[3]), .o_cout(cout21[3]));
pu pu21_4 (.i_a(result20[3]), .i_b(~i_divisor[4]), .i_cin(cout21[3]), .i_carry_output(quotient[10]),
		.o_result(result21[4]), .o_cout(cout21[4]));
pu pu21_5 (.i_a(result20[4]), .i_b(~i_divisor[5]), .i_cin(cout21[4]), .i_carry_output(quotient[10]),
		.o_result(result21[5]), .o_cout(cout21[5]));
pu pu21_6 (.i_a(result20[5]), .i_b(~i_divisor[6]), .i_cin(cout21[5]), .i_carry_output(quotient[10]),
		.o_result(result21[6]), .o_cout(cout21[6]));
pu pu21_7 (.i_a(result20[6]), .i_b(~i_divisor[7]), .i_cin(cout21[6]), .i_carry_output(quotient[10]),
		.o_result(result21[7]), .o_cout(cout21[7]));
pu pu21_8 (.i_a(result20[7]), .i_b(~i_divisor[8]), .i_cin(cout21[7]), .i_carry_output(quotient[10]),
		.o_result(result21[8]), .o_cout(cout21[8]));
pu pu21_9 (.i_a(result20[8]), .i_b(~i_divisor[9]), .i_cin(cout21[8]), .i_carry_output(quotient[10]),
		.o_result(result21[9]), .o_cout(cout21[9]));
pu pu21_10 (.i_a(result20[9]), .i_b(~i_divisor[10]), .i_cin(cout21[9]), .i_carry_output(quotient[10]),
		.o_result(result21[10]), .o_cout(cout21[10]));
pu pu21_11 (.i_a(result20[10]), .i_b(~i_divisor[11]), .i_cin(cout21[10]), .i_carry_output(quotient[10]),
		.o_result(result21[11]), .o_cout(cout21[11]));
pu pu21_12 (.i_a(result20[11]), .i_b(~i_divisor[12]), .i_cin(cout21[11]), .i_carry_output(quotient[10]),
		.o_result(result21[12]), .o_cout(cout21[12]));
pu pu21_13 (.i_a(result20[12]), .i_b(~i_divisor[13]), .i_cin(cout21[12]), .i_carry_output(quotient[10]),
		.o_result(result21[13]), .o_cout(cout21[13]));
pu pu21_14 (.i_a(result20[13]), .i_b(~i_divisor[14]), .i_cin(cout21[13]), .i_carry_output(quotient[10]),
		.o_result(result21[14]), .o_cout(cout21[14]));
pu pu21_15 (.i_a(result20[14]), .i_b(~i_divisor[15]), .i_cin(cout21[14]), .i_carry_output(quotient[10]),
		.o_result(result21[15]), .o_cout(cout21[15]));
pu pu21_16 (.i_a(result20[15]), .i_b(~i_divisor[16]), .i_cin(cout21[15]), .i_carry_output(quotient[10]),
		.o_result(result21[16]), .o_cout(cout21[16]));
pu pu21_17 (.i_a(result20[16]), .i_b(~i_divisor[17]), .i_cin(cout21[16]), .i_carry_output(quotient[10]),
		.o_result(result21[17]), .o_cout(cout21[17]));
pu pu21_18 (.i_a(result20[17]), .i_b(~i_divisor[18]), .i_cin(cout21[17]), .i_carry_output(quotient[10]),
		.o_result(result21[18]), .o_cout(cout21[18]));
pu pu21_19 (.i_a(result20[18]), .i_b(~i_divisor[19]), .i_cin(cout21[18]), .i_carry_output(quotient[10]),
		.o_result(result21[19]), .o_cout(cout21[19]));
pu pu21_20 (.i_a(result20[19]), .i_b(~i_divisor[20]), .i_cin(cout21[19]), .i_carry_output(quotient[10]),
		.o_result(result21[20]), .o_cout(cout21[20]));
pu pu21_21 (.i_a(result20[20]), .i_b(~i_divisor[21]), .i_cin(cout21[20]), .i_carry_output(quotient[10]),
		.o_result(result21[21]), .o_cout(cout21[21]));
pu pu21_22 (.i_a(result20[21]), .i_b(~i_divisor[22]), .i_cin(cout21[21]), .i_carry_output(quotient[10]),
		.o_result(result21[22]), .o_cout(cout21[22]));
pu pu21_23 (.i_a(result20[22]), .i_b(~i_divisor[23]), .i_cin(cout21[22]), .i_carry_output(quotient[10]),
		.o_result(result21[23]), .o_cout(cout21[23]));
pu pu21_24 (.i_a(result20[23]), .i_b(~i_divisor[24]), .i_cin(cout21[23]), .i_carry_output(quotient[10]),
		.o_result(result21[24]), .o_cout(cout21[24]));
pu pu21_25 (.i_a(result20[24]), .i_b(~i_divisor[25]), .i_cin(cout21[24]), .i_carry_output(quotient[10]),
		.o_result(result21[25]), .o_cout(cout21[25]));
pu pu21_26 (.i_a(result20[25]), .i_b(~i_divisor[26]), .i_cin(cout21[25]), .i_carry_output(quotient[10]),
		.o_result(result21[26]), .o_cout(cout21[26]));
pu pu21_27 (.i_a(result20[26]), .i_b(~i_divisor[27]), .i_cin(cout21[26]), .i_carry_output(quotient[10]),
		.o_result(result21[27]), .o_cout(cout21[27]));
pu pu21_28 (.i_a(result20[27]), .i_b(~i_divisor[28]), .i_cin(cout21[27]), .i_carry_output(quotient[10]),
		.o_result(result21[28]), .o_cout(cout21[28]));
pu pu21_29 (.i_a(result20[28]), .i_b(~i_divisor[29]), .i_cin(cout21[28]), .i_carry_output(quotient[10]),
		.o_result(result21[29]), .o_cout(cout21[29]));
pu pu21_30 (.i_a(result20[29]), .i_b(~i_divisor[30]), .i_cin(cout21[29]), .i_carry_output(quotient[10]),
		.o_result(result21[30]), .o_cout(cout21[30]));
pu pu21_31 (.i_a(result20[30]), .i_b(~i_divisor[31]), .i_cin(cout21[30]), .i_carry_output(quotient[10]),
		.o_cout(quotient[10]));

// Row 22
pu pu22_0 (.i_a(i_dividend[9]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[9]),
         .o_result(result22[0]), .o_cout(cout22[0]));
pu pu22_1 (.i_a(result21[0]), .i_b(~i_divisor[1]), .i_cin(cout22[0]), .i_carry_output(quotient[9]),
		.o_result(result22[1]), .o_cout(cout22[1]));
pu pu22_2 (.i_a(result21[1]), .i_b(~i_divisor[2]), .i_cin(cout22[1]), .i_carry_output(quotient[9]),
		.o_result(result22[2]), .o_cout(cout22[2]));
pu pu22_3 (.i_a(result21[2]), .i_b(~i_divisor[3]), .i_cin(cout22[2]), .i_carry_output(quotient[9]),
		.o_result(result22[3]), .o_cout(cout22[3]));
pu pu22_4 (.i_a(result21[3]), .i_b(~i_divisor[4]), .i_cin(cout22[3]), .i_carry_output(quotient[9]),
		.o_result(result22[4]), .o_cout(cout22[4]));
pu pu22_5 (.i_a(result21[4]), .i_b(~i_divisor[5]), .i_cin(cout22[4]), .i_carry_output(quotient[9]),
		.o_result(result22[5]), .o_cout(cout22[5]));
pu pu22_6 (.i_a(result21[5]), .i_b(~i_divisor[6]), .i_cin(cout22[5]), .i_carry_output(quotient[9]),
		.o_result(result22[6]), .o_cout(cout22[6]));
pu pu22_7 (.i_a(result21[6]), .i_b(~i_divisor[7]), .i_cin(cout22[6]), .i_carry_output(quotient[9]),
		.o_result(result22[7]), .o_cout(cout22[7]));
pu pu22_8 (.i_a(result21[7]), .i_b(~i_divisor[8]), .i_cin(cout22[7]), .i_carry_output(quotient[9]),
		.o_result(result22[8]), .o_cout(cout22[8]));
pu pu22_9 (.i_a(result21[8]), .i_b(~i_divisor[9]), .i_cin(cout22[8]), .i_carry_output(quotient[9]),
		.o_result(result22[9]), .o_cout(cout22[9]));
pu pu22_10 (.i_a(result21[9]), .i_b(~i_divisor[10]), .i_cin(cout22[9]), .i_carry_output(quotient[9]),
		.o_result(result22[10]), .o_cout(cout22[10]));
pu pu22_11 (.i_a(result21[10]), .i_b(~i_divisor[11]), .i_cin(cout22[10]), .i_carry_output(quotient[9]),
		.o_result(result22[11]), .o_cout(cout22[11]));
pu pu22_12 (.i_a(result21[11]), .i_b(~i_divisor[12]), .i_cin(cout22[11]), .i_carry_output(quotient[9]),
		.o_result(result22[12]), .o_cout(cout22[12]));
pu pu22_13 (.i_a(result21[12]), .i_b(~i_divisor[13]), .i_cin(cout22[12]), .i_carry_output(quotient[9]),
		.o_result(result22[13]), .o_cout(cout22[13]));
pu pu22_14 (.i_a(result21[13]), .i_b(~i_divisor[14]), .i_cin(cout22[13]), .i_carry_output(quotient[9]),
		.o_result(result22[14]), .o_cout(cout22[14]));
pu pu22_15 (.i_a(result21[14]), .i_b(~i_divisor[15]), .i_cin(cout22[14]), .i_carry_output(quotient[9]),
		.o_result(result22[15]), .o_cout(cout22[15]));
pu pu22_16 (.i_a(result21[15]), .i_b(~i_divisor[16]), .i_cin(cout22[15]), .i_carry_output(quotient[9]),
		.o_result(result22[16]), .o_cout(cout22[16]));
pu pu22_17 (.i_a(result21[16]), .i_b(~i_divisor[17]), .i_cin(cout22[16]), .i_carry_output(quotient[9]),
		.o_result(result22[17]), .o_cout(cout22[17]));
pu pu22_18 (.i_a(result21[17]), .i_b(~i_divisor[18]), .i_cin(cout22[17]), .i_carry_output(quotient[9]),
		.o_result(result22[18]), .o_cout(cout22[18]));
pu pu22_19 (.i_a(result21[18]), .i_b(~i_divisor[19]), .i_cin(cout22[18]), .i_carry_output(quotient[9]),
		.o_result(result22[19]), .o_cout(cout22[19]));
pu pu22_20 (.i_a(result21[19]), .i_b(~i_divisor[20]), .i_cin(cout22[19]), .i_carry_output(quotient[9]),
		.o_result(result22[20]), .o_cout(cout22[20]));
pu pu22_21 (.i_a(result21[20]), .i_b(~i_divisor[21]), .i_cin(cout22[20]), .i_carry_output(quotient[9]),
		.o_result(result22[21]), .o_cout(cout22[21]));
pu pu22_22 (.i_a(result21[21]), .i_b(~i_divisor[22]), .i_cin(cout22[21]), .i_carry_output(quotient[9]),
		.o_result(result22[22]), .o_cout(cout22[22]));
pu pu22_23 (.i_a(result21[22]), .i_b(~i_divisor[23]), .i_cin(cout22[22]), .i_carry_output(quotient[9]),
		.o_result(result22[23]), .o_cout(cout22[23]));
pu pu22_24 (.i_a(result21[23]), .i_b(~i_divisor[24]), .i_cin(cout22[23]), .i_carry_output(quotient[9]),
		.o_result(result22[24]), .o_cout(cout22[24]));
pu pu22_25 (.i_a(result21[24]), .i_b(~i_divisor[25]), .i_cin(cout22[24]), .i_carry_output(quotient[9]),
		.o_result(result22[25]), .o_cout(cout22[25]));
pu pu22_26 (.i_a(result21[25]), .i_b(~i_divisor[26]), .i_cin(cout22[25]), .i_carry_output(quotient[9]),
		.o_result(result22[26]), .o_cout(cout22[26]));
pu pu22_27 (.i_a(result21[26]), .i_b(~i_divisor[27]), .i_cin(cout22[26]), .i_carry_output(quotient[9]),
		.o_result(result22[27]), .o_cout(cout22[27]));
pu pu22_28 (.i_a(result21[27]), .i_b(~i_divisor[28]), .i_cin(cout22[27]), .i_carry_output(quotient[9]),
		.o_result(result22[28]), .o_cout(cout22[28]));
pu pu22_29 (.i_a(result21[28]), .i_b(~i_divisor[29]), .i_cin(cout22[28]), .i_carry_output(quotient[9]),
		.o_result(result22[29]), .o_cout(cout22[29]));
pu pu22_30 (.i_a(result21[29]), .i_b(~i_divisor[30]), .i_cin(cout22[29]), .i_carry_output(quotient[9]),
		.o_result(result22[30]), .o_cout(cout22[30]));
pu pu22_31 (.i_a(result21[30]), .i_b(~i_divisor[31]), .i_cin(cout22[30]), .i_carry_output(quotient[9]),
		.o_cout(quotient[9]));

// Row 23
pu pu23_0 (.i_a(i_dividend[8]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[8]),
         .o_result(result23[0]), .o_cout(cout23[0]));
pu pu23_1 (.i_a(result22[0]), .i_b(~i_divisor[1]), .i_cin(cout23[0]), .i_carry_output(quotient[8]),
		.o_result(result23[1]), .o_cout(cout23[1]));
pu pu23_2 (.i_a(result22[1]), .i_b(~i_divisor[2]), .i_cin(cout23[1]), .i_carry_output(quotient[8]),
		.o_result(result23[2]), .o_cout(cout23[2]));
pu pu23_3 (.i_a(result22[2]), .i_b(~i_divisor[3]), .i_cin(cout23[2]), .i_carry_output(quotient[8]),
		.o_result(result23[3]), .o_cout(cout23[3]));
pu pu23_4 (.i_a(result22[3]), .i_b(~i_divisor[4]), .i_cin(cout23[3]), .i_carry_output(quotient[8]),
		.o_result(result23[4]), .o_cout(cout23[4]));
pu pu23_5 (.i_a(result22[4]), .i_b(~i_divisor[5]), .i_cin(cout23[4]), .i_carry_output(quotient[8]),
		.o_result(result23[5]), .o_cout(cout23[5]));
pu pu23_6 (.i_a(result22[5]), .i_b(~i_divisor[6]), .i_cin(cout23[5]), .i_carry_output(quotient[8]),
		.o_result(result23[6]), .o_cout(cout23[6]));
pu pu23_7 (.i_a(result22[6]), .i_b(~i_divisor[7]), .i_cin(cout23[6]), .i_carry_output(quotient[8]),
		.o_result(result23[7]), .o_cout(cout23[7]));
pu pu23_8 (.i_a(result22[7]), .i_b(~i_divisor[8]), .i_cin(cout23[7]), .i_carry_output(quotient[8]),
		.o_result(result23[8]), .o_cout(cout23[8]));
pu pu23_9 (.i_a(result22[8]), .i_b(~i_divisor[9]), .i_cin(cout23[8]), .i_carry_output(quotient[8]),
		.o_result(result23[9]), .o_cout(cout23[9]));
pu pu23_10 (.i_a(result22[9]), .i_b(~i_divisor[10]), .i_cin(cout23[9]), .i_carry_output(quotient[8]),
		.o_result(result23[10]), .o_cout(cout23[10]));
pu pu23_11 (.i_a(result22[10]), .i_b(~i_divisor[11]), .i_cin(cout23[10]), .i_carry_output(quotient[8]),
		.o_result(result23[11]), .o_cout(cout23[11]));
pu pu23_12 (.i_a(result22[11]), .i_b(~i_divisor[12]), .i_cin(cout23[11]), .i_carry_output(quotient[8]),
		.o_result(result23[12]), .o_cout(cout23[12]));
pu pu23_13 (.i_a(result22[12]), .i_b(~i_divisor[13]), .i_cin(cout23[12]), .i_carry_output(quotient[8]),
		.o_result(result23[13]), .o_cout(cout23[13]));
pu pu23_14 (.i_a(result22[13]), .i_b(~i_divisor[14]), .i_cin(cout23[13]), .i_carry_output(quotient[8]),
		.o_result(result23[14]), .o_cout(cout23[14]));
pu pu23_15 (.i_a(result22[14]), .i_b(~i_divisor[15]), .i_cin(cout23[14]), .i_carry_output(quotient[8]),
		.o_result(result23[15]), .o_cout(cout23[15]));
pu pu23_16 (.i_a(result22[15]), .i_b(~i_divisor[16]), .i_cin(cout23[15]), .i_carry_output(quotient[8]),
		.o_result(result23[16]), .o_cout(cout23[16]));
pu pu23_17 (.i_a(result22[16]), .i_b(~i_divisor[17]), .i_cin(cout23[16]), .i_carry_output(quotient[8]),
		.o_result(result23[17]), .o_cout(cout23[17]));
pu pu23_18 (.i_a(result22[17]), .i_b(~i_divisor[18]), .i_cin(cout23[17]), .i_carry_output(quotient[8]),
		.o_result(result23[18]), .o_cout(cout23[18]));
pu pu23_19 (.i_a(result22[18]), .i_b(~i_divisor[19]), .i_cin(cout23[18]), .i_carry_output(quotient[8]),
		.o_result(result23[19]), .o_cout(cout23[19]));
pu pu23_20 (.i_a(result22[19]), .i_b(~i_divisor[20]), .i_cin(cout23[19]), .i_carry_output(quotient[8]),
		.o_result(result23[20]), .o_cout(cout23[20]));
pu pu23_21 (.i_a(result22[20]), .i_b(~i_divisor[21]), .i_cin(cout23[20]), .i_carry_output(quotient[8]),
		.o_result(result23[21]), .o_cout(cout23[21]));
pu pu23_22 (.i_a(result22[21]), .i_b(~i_divisor[22]), .i_cin(cout23[21]), .i_carry_output(quotient[8]),
		.o_result(result23[22]), .o_cout(cout23[22]));
pu pu23_23 (.i_a(result22[22]), .i_b(~i_divisor[23]), .i_cin(cout23[22]), .i_carry_output(quotient[8]),
		.o_result(result23[23]), .o_cout(cout23[23]));
pu pu23_24 (.i_a(result22[23]), .i_b(~i_divisor[24]), .i_cin(cout23[23]), .i_carry_output(quotient[8]),
		.o_result(result23[24]), .o_cout(cout23[24]));
pu pu23_25 (.i_a(result22[24]), .i_b(~i_divisor[25]), .i_cin(cout23[24]), .i_carry_output(quotient[8]),
		.o_result(result23[25]), .o_cout(cout23[25]));
pu pu23_26 (.i_a(result22[25]), .i_b(~i_divisor[26]), .i_cin(cout23[25]), .i_carry_output(quotient[8]),
		.o_result(result23[26]), .o_cout(cout23[26]));
pu pu23_27 (.i_a(result22[26]), .i_b(~i_divisor[27]), .i_cin(cout23[26]), .i_carry_output(quotient[8]),
		.o_result(result23[27]), .o_cout(cout23[27]));
pu pu23_28 (.i_a(result22[27]), .i_b(~i_divisor[28]), .i_cin(cout23[27]), .i_carry_output(quotient[8]),
		.o_result(result23[28]), .o_cout(cout23[28]));
pu pu23_29 (.i_a(result22[28]), .i_b(~i_divisor[29]), .i_cin(cout23[28]), .i_carry_output(quotient[8]),
		.o_result(result23[29]), .o_cout(cout23[29]));
pu pu23_30 (.i_a(result22[29]), .i_b(~i_divisor[30]), .i_cin(cout23[29]), .i_carry_output(quotient[8]),
		.o_result(result23[30]), .o_cout(cout23[30]));
pu pu23_31 (.i_a(result22[30]), .i_b(~i_divisor[31]), .i_cin(cout23[30]), .i_carry_output(quotient[8]),
		.o_cout(quotient[8]));

// Row 24
pu pu24_0 (.i_a(i_dividend[7]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[7]),
         .o_result(result24[0]), .o_cout(cout24[0]));	
pu pu24_1 (.i_a(result23[0]), .i_b(~i_divisor[1]), .i_cin(cout24[0]), .i_carry_output(quotient[7]),
		.o_result(result24[1]), .o_cout(cout24[1]));
pu pu24_2 (.i_a(result23[1]), .i_b(~i_divisor[2]), .i_cin(cout24[1]), .i_carry_output(quotient[7]),
		.o_result(result24[2]), .o_cout(cout24[2]));
pu pu24_3 (.i_a(result23[2]), .i_b(~i_divisor[3]), .i_cin(cout24[2]), .i_carry_output(quotient[7]),
		.o_result(result24[3]), .o_cout(cout24[3]));
pu pu24_4 (.i_a(result23[3]), .i_b(~i_divisor[4]), .i_cin(cout24[3]), .i_carry_output(quotient[7]),
		.o_result(result24[4]), .o_cout(cout24[4]));
pu pu24_5 (.i_a(result23[4]), .i_b(~i_divisor[5]), .i_cin(cout24[4]), .i_carry_output(quotient[7]),
		.o_result(result24[5]), .o_cout(cout24[5]));
pu pu24_6 (.i_a(result23[5]), .i_b(~i_divisor[6]), .i_cin(cout24[5]), .i_carry_output(quotient[7]),
		.o_result(result24[6]), .o_cout(cout24[6]));
pu pu24_7 (.i_a(result23[6]), .i_b(~i_divisor[7]), .i_cin(cout24[6]), .i_carry_output(quotient[7]),
		.o_result(result24[7]), .o_cout(cout24[7]));
pu pu24_8 (.i_a(result23[7]), .i_b(~i_divisor[8]), .i_cin(cout24[7]), .i_carry_output(quotient[7]),
		.o_result(result24[8]), .o_cout(cout24[8]));
pu pu24_9 (.i_a(result23[8]), .i_b(~i_divisor[9]), .i_cin(cout24[8]), .i_carry_output(quotient[7]),
		.o_result(result24[9]), .o_cout(cout24[9]));
pu pu24_10 (.i_a(result23[9]), .i_b(~i_divisor[10]), .i_cin(cout24[9]), .i_carry_output(quotient[7]),
		.o_result(result24[10]), .o_cout(cout24[10]));
pu pu24_11 (.i_a(result23[10]), .i_b(~i_divisor[11]), .i_cin(cout24[10]), .i_carry_output(quotient[7]),
		.o_result(result24[11]), .o_cout(cout24[11]));
pu pu24_12 (.i_a(result23[11]), .i_b(~i_divisor[12]), .i_cin(cout24[11]), .i_carry_output(quotient[7]),
		.o_result(result24[12]), .o_cout(cout24[12]));
pu pu24_13 (.i_a(result23[12]), .i_b(~i_divisor[13]), .i_cin(cout24[12]), .i_carry_output(quotient[7]),
		.o_result(result24[13]), .o_cout(cout24[13]));
pu pu24_14 (.i_a(result23[13]), .i_b(~i_divisor[14]), .i_cin(cout24[13]), .i_carry_output(quotient[7]),
		.o_result(result24[14]), .o_cout(cout24[14]));
pu pu24_15 (.i_a(result23[14]), .i_b(~i_divisor[15]), .i_cin(cout24[14]), .i_carry_output(quotient[7]),
		.o_result(result24[15]), .o_cout(cout24[15]));
pu pu24_16 (.i_a(result23[15]), .i_b(~i_divisor[16]), .i_cin(cout24[15]), .i_carry_output(quotient[7]),
		.o_result(result24[16]), .o_cout(cout24[16]));
pu pu24_17 (.i_a(result23[16]), .i_b(~i_divisor[17]), .i_cin(cout24[16]), .i_carry_output(quotient[7]),
		.o_result(result24[17]), .o_cout(cout24[17]));
pu pu24_18 (.i_a(result23[17]), .i_b(~i_divisor[18]), .i_cin(cout24[17]), .i_carry_output(quotient[7]),
		.o_result(result24[18]), .o_cout(cout24[18]));
pu pu24_19 (.i_a(result23[18]), .i_b(~i_divisor[19]), .i_cin(cout24[18]), .i_carry_output(quotient[7]),
		.o_result(result24[19]), .o_cout(cout24[19]));
pu pu24_20 (.i_a(result23[19]), .i_b(~i_divisor[20]), .i_cin(cout24[19]), .i_carry_output(quotient[7]),
		.o_result(result24[20]), .o_cout(cout24[20]));
pu pu24_21 (.i_a(result23[20]), .i_b(~i_divisor[21]), .i_cin(cout24[20]), .i_carry_output(quotient[7]),
		.o_result(result24[21]), .o_cout(cout24[21]));
pu pu24_22 (.i_a(result23[21]), .i_b(~i_divisor[22]), .i_cin(cout24[21]), .i_carry_output(quotient[7]),
		.o_result(result24[22]), .o_cout(cout24[22]));
pu pu24_23 (.i_a(result23[22]), .i_b(~i_divisor[23]), .i_cin(cout24[22]), .i_carry_output(quotient[7]),
		.o_result(result24[23]), .o_cout(cout24[23]));
pu pu24_24 (.i_a(result23[23]), .i_b(~i_divisor[24]), .i_cin(cout24[23]), .i_carry_output(quotient[7]),
		.o_result(result24[24]), .o_cout(cout24[24]));
pu pu24_25 (.i_a(result23[24]), .i_b(~i_divisor[25]), .i_cin(cout24[24]), .i_carry_output(quotient[7]),
		.o_result(result24[25]), .o_cout(cout24[25]));
pu pu24_26 (.i_a(result23[25]), .i_b(~i_divisor[26]), .i_cin(cout24[25]), .i_carry_output(quotient[7]),
		.o_result(result24[26]), .o_cout(cout24[26]));
pu pu24_27 (.i_a(result23[26]), .i_b(~i_divisor[27]), .i_cin(cout24[26]), .i_carry_output(quotient[7]),
		.o_result(result24[27]), .o_cout(cout24[27]));
pu pu24_28 (.i_a(result23[27]), .i_b(~i_divisor[28]), .i_cin(cout24[27]), .i_carry_output(quotient[7]),
		.o_result(result24[28]), .o_cout(cout24[28]));
pu pu24_29 (.i_a(result23[28]), .i_b(~i_divisor[29]), .i_cin(cout24[28]), .i_carry_output(quotient[7]),
		.o_result(result24[29]), .o_cout(cout24[29]));
pu pu24_30 (.i_a(result23[29]), .i_b(~i_divisor[30]), .i_cin(cout24[29]), .i_carry_output(quotient[7]),
		.o_result(result24[30]), .o_cout(cout24[30]));
pu pu24_31 (.i_a(result23[30]), .i_b(~i_divisor[31]), .i_cin(cout24[30]), .i_carry_output(quotient[7]),
		.o_cout(quotient[7]));

// Row 25
pu pu25_0 (.i_a(i_dividend[6]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[6]),
         .o_result(result25[0]), .o_cout(cout25[0]));	
pu pu25_1 (.i_a(result24[0]), .i_b(~i_divisor[1]), .i_cin(cout25[0]), .i_carry_output(quotient[6]),
		.o_result(result25[1]), .o_cout(cout25[1]));
pu pu25_2 (.i_a(result24[1]), .i_b(~i_divisor[2]), .i_cin(cout25[1]), .i_carry_output(quotient[6]),
		.o_result(result25[2]), .o_cout(cout25[2]));
pu pu25_3 (.i_a(result24[2]), .i_b(~i_divisor[3]), .i_cin(cout25[2]), .i_carry_output(quotient[6]),
		.o_result(result25[3]), .o_cout(cout25[3]));
pu pu25_4 (.i_a(result24[3]), .i_b(~i_divisor[4]), .i_cin(cout25[3]), .i_carry_output(quotient[6]),
		.o_result(result25[4]), .o_cout(cout25[4]));
pu pu25_5 (.i_a(result24[4]), .i_b(~i_divisor[5]), .i_cin(cout25[4]), .i_carry_output(quotient[6]),
		.o_result(result25[5]), .o_cout(cout25[5]));
pu pu25_6 (.i_a(result24[5]), .i_b(~i_divisor[6]), .i_cin(cout25[5]), .i_carry_output(quotient[6]),
		.o_result(result25[6]), .o_cout(cout25[6]));
pu pu25_7 (.i_a(result24[6]), .i_b(~i_divisor[7]), .i_cin(cout25[6]), .i_carry_output(quotient[6]),
		.o_result(result25[7]), .o_cout(cout25[7]));
pu pu25_8 (.i_a(result24[7]), .i_b(~i_divisor[8]), .i_cin(cout25[7]), .i_carry_output(quotient[6]),
		.o_result(result25[8]), .o_cout(cout25[8]));
pu pu25_9 (.i_a(result24[8]), .i_b(~i_divisor[9]), .i_cin(cout25[8]), .i_carry_output(quotient[6]),
		.o_result(result25[9]), .o_cout(cout25[9]));
pu pu25_10 (.i_a(result24[9]), .i_b(~i_divisor[10]), .i_cin(cout25[9]), .i_carry_output(quotient[6]),
		.o_result(result25[10]), .o_cout(cout25[10]));
pu pu25_11 (.i_a(result24[10]), .i_b(~i_divisor[11]), .i_cin(cout25[10]), .i_carry_output(quotient[6]),
		.o_result(result25[11]), .o_cout(cout25[11]));
pu pu25_12 (.i_a(result24[11]), .i_b(~i_divisor[12]), .i_cin(cout25[11]), .i_carry_output(quotient[6]),
		.o_result(result25[12]), .o_cout(cout25[12]));
pu pu25_13 (.i_a(result24[12]), .i_b(~i_divisor[13]), .i_cin(cout25[12]), .i_carry_output(quotient[6]),
		.o_result(result25[13]), .o_cout(cout25[13]));
pu pu25_14 (.i_a(result24[13]), .i_b(~i_divisor[14]), .i_cin(cout25[13]), .i_carry_output(quotient[6]),
		.o_result(result25[14]), .o_cout(cout25[14]));
pu pu25_15 (.i_a(result24[14]), .i_b(~i_divisor[15]), .i_cin(cout25[14]), .i_carry_output(quotient[6]),
		.o_result(result25[15]), .o_cout(cout25[15]));
pu pu25_16 (.i_a(result24[15]), .i_b(~i_divisor[16]), .i_cin(cout25[15]), .i_carry_output(quotient[6]),
		.o_result(result25[16]), .o_cout(cout25[16]));
pu pu25_17 (.i_a(result24[16]), .i_b(~i_divisor[17]), .i_cin(cout25[16]), .i_carry_output(quotient[6]),
		.o_result(result25[17]), .o_cout(cout25[17]));
pu pu25_18 (.i_a(result24[17]), .i_b(~i_divisor[18]), .i_cin(cout25[17]), .i_carry_output(quotient[6]),
		.o_result(result25[18]), .o_cout(cout25[18]));
pu pu25_19 (.i_a(result24[18]), .i_b(~i_divisor[19]), .i_cin(cout25[18]), .i_carry_output(quotient[6]),
		.o_result(result25[19]), .o_cout(cout25[19]));
pu pu25_20 (.i_a(result24[19]), .i_b(~i_divisor[20]), .i_cin(cout25[19]), .i_carry_output(quotient[6]),
		.o_result(result25[20]), .o_cout(cout25[20]));
pu pu25_21 (.i_a(result24[20]), .i_b(~i_divisor[21]), .i_cin(cout25[20]), .i_carry_output(quotient[6]),
		.o_result(result25[21]), .o_cout(cout25[21]));
pu pu25_22 (.i_a(result24[21]), .i_b(~i_divisor[22]), .i_cin(cout25[21]), .i_carry_output(quotient[6]),
		.o_result(result25[22]), .o_cout(cout25[22]));
pu pu25_23 (.i_a(result24[22]), .i_b(~i_divisor[23]), .i_cin(cout25[22]), .i_carry_output(quotient[6]),
		.o_result(result25[23]), .o_cout(cout25[23]));
pu pu25_24 (.i_a(result24[23]), .i_b(~i_divisor[24]), .i_cin(cout25[23]), .i_carry_output(quotient[6]),
		.o_result(result25[24]), .o_cout(cout25[24]));
pu pu25_25 (.i_a(result24[24]), .i_b(~i_divisor[25]), .i_cin(cout25[24]), .i_carry_output(quotient[6]),
		.o_result(result25[25]), .o_cout(cout25[25]));
pu pu25_26 (.i_a(result24[25]), .i_b(~i_divisor[26]), .i_cin(cout25[25]), .i_carry_output(quotient[6]),
		.o_result(result25[26]), .o_cout(cout25[26]));
pu pu25_27 (.i_a(result24[26]), .i_b(~i_divisor[27]), .i_cin(cout25[26]), .i_carry_output(quotient[6]),
		.o_result(result25[27]), .o_cout(cout25[27]));
pu pu25_28 (.i_a(result24[27]), .i_b(~i_divisor[28]), .i_cin(cout25[27]), .i_carry_output(quotient[6]),
		.o_result(result25[28]), .o_cout(cout25[28]));
pu pu25_29 (.i_a(result24[28]), .i_b(~i_divisor[29]), .i_cin(cout25[28]), .i_carry_output(quotient[6]),
		.o_result(result25[29]), .o_cout(cout25[29]));
pu pu25_30 (.i_a(result24[29]), .i_b(~i_divisor[30]), .i_cin(cout25[29]), .i_carry_output(quotient[6]),
		.o_result(result25[30]), .o_cout(cout25[30]));
pu pu25_31 (.i_a(result24[30]), .i_b(~i_divisor[31]), .i_cin(cout25[30]), .i_carry_output(quotient[6]),
		.o_cout(quotient[6]));

// Row 26
pu pu26_0 (.i_a(i_dividend[5]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[5]),
         .o_result(result26[0]), .o_cout(cout26[0]));	
pu pu26_1 (.i_a(result25[0]), .i_b(~i_divisor[1]), .i_cin(cout26[0]), .i_carry_output(quotient[5]),
		.o_result(result26[1]), .o_cout(cout26[1]));
pu pu26_2 (.i_a(result25[1]), .i_b(~i_divisor[2]), .i_cin(cout26[1]), .i_carry_output(quotient[5]),
		.o_result(result26[2]), .o_cout(cout26[2]));
pu pu26_3 (.i_a(result25[2]), .i_b(~i_divisor[3]), .i_cin(cout26[2]), .i_carry_output(quotient[5]),
		.o_result(result26[3]), .o_cout(cout26[3]));
pu pu26_4 (.i_a(result25[3]), .i_b(~i_divisor[4]), .i_cin(cout26[3]), .i_carry_output(quotient[5]),
		.o_result(result26[4]), .o_cout(cout26[4]));
pu pu26_5 (.i_a(result25[4]), .i_b(~i_divisor[5]), .i_cin(cout26[4]), .i_carry_output(quotient[5]),
		.o_result(result26[5]), .o_cout(cout26[5]));
pu pu26_6 (.i_a(result25[5]), .i_b(~i_divisor[6]), .i_cin(cout26[5]), .i_carry_output(quotient[5]),
		.o_result(result26[6]), .o_cout(cout26[6]));
pu pu26_7 (.i_a(result25[6]), .i_b(~i_divisor[7]), .i_cin(cout26[6]), .i_carry_output(quotient[5]),
		.o_result(result26[7]), .o_cout(cout26[7]));
pu pu26_8 (.i_a(result25[7]), .i_b(~i_divisor[8]), .i_cin(cout26[7]), .i_carry_output(quotient[5]),
		.o_result(result26[8]), .o_cout(cout26[8]));
pu pu26_9 (.i_a(result25[8]), .i_b(~i_divisor[9]), .i_cin(cout26[8]), .i_carry_output(quotient[5]),
		.o_result(result26[9]), .o_cout(cout26[9]));
pu pu26_10 (.i_a(result25[9]), .i_b(~i_divisor[10]), .i_cin(cout26[9]), .i_carry_output(quotient[5]),
		.o_result(result26[10]), .o_cout(cout26[10]));
pu pu26_11 (.i_a(result25[10]), .i_b(~i_divisor[11]), .i_cin(cout26[10]), .i_carry_output(quotient[5]),
		.o_result(result26[11]), .o_cout(cout26[11]));
pu pu26_12 (.i_a(result25[11]), .i_b(~i_divisor[12]), .i_cin(cout26[11]), .i_carry_output(quotient[5]),
		.o_result(result26[12]), .o_cout(cout26[12]));
pu pu26_13 (.i_a(result25[12]), .i_b(~i_divisor[13]), .i_cin(cout26[12]), .i_carry_output(quotient[5]),
		.o_result(result26[13]), .o_cout(cout26[13]));
pu pu26_14 (.i_a(result25[13]), .i_b(~i_divisor[14]), .i_cin(cout26[13]), .i_carry_output(quotient[5]),
		.o_result(result26[14]), .o_cout(cout26[14]));
pu pu26_15 (.i_a(result25[14]), .i_b(~i_divisor[15]), .i_cin(cout26[14]), .i_carry_output(quotient[5]),
		.o_result(result26[15]), .o_cout(cout26[15]));
pu pu26_16 (.i_a(result25[15]), .i_b(~i_divisor[16]), .i_cin(cout26[15]), .i_carry_output(quotient[5]),
		.o_result(result26[16]), .o_cout(cout26[16]));
pu pu26_17 (.i_a(result25[16]), .i_b(~i_divisor[17]), .i_cin(cout26[16]), .i_carry_output(quotient[5]),
		.o_result(result26[17]), .o_cout(cout26[17]));
pu pu26_18 (.i_a(result25[17]), .i_b(~i_divisor[18]), .i_cin(cout26[17]), .i_carry_output(quotient[5]),
		.o_result(result26[18]), .o_cout(cout26[18]));
pu pu26_19 (.i_a(result25[18]), .i_b(~i_divisor[19]), .i_cin(cout26[18]), .i_carry_output(quotient[5]),
		.o_result(result26[19]), .o_cout(cout26[19]));
pu pu26_20 (.i_a(result25[19]), .i_b(~i_divisor[20]), .i_cin(cout26[19]), .i_carry_output(quotient[5]),
		.o_result(result26[20]), .o_cout(cout26[20]));
pu pu26_21 (.i_a(result25[20]), .i_b(~i_divisor[21]), .i_cin(cout26[20]), .i_carry_output(quotient[5]),
		.o_result(result26[21]), .o_cout(cout26[21]));
pu pu26_22 (.i_a(result25[21]), .i_b(~i_divisor[22]), .i_cin(cout26[21]), .i_carry_output(quotient[5]),
		.o_result(result26[22]), .o_cout(cout26[22]));
pu pu26_23 (.i_a(result25[22]), .i_b(~i_divisor[23]), .i_cin(cout26[22]), .i_carry_output(quotient[5]),
		.o_result(result26[23]), .o_cout(cout26[23]));
pu pu26_24 (.i_a(result25[23]), .i_b(~i_divisor[24]), .i_cin(cout26[23]), .i_carry_output(quotient[5]),
		.o_result(result26[24]), .o_cout(cout26[24]));
pu pu26_25 (.i_a(result25[24]), .i_b(~i_divisor[25]), .i_cin(cout26[24]), .i_carry_output(quotient[5]),
		.o_result(result26[25]), .o_cout(cout26[25]));
pu pu26_26 (.i_a(result25[25]), .i_b(~i_divisor[26]), .i_cin(cout26[25]), .i_carry_output(quotient[5]),
		.o_result(result26[26]), .o_cout(cout26[26]));
pu pu26_27 (.i_a(result25[26]), .i_b(~i_divisor[27]), .i_cin(cout26[26]), .i_carry_output(quotient[5]),
		.o_result(result26[27]), .o_cout(cout26[27]));
pu pu26_28 (.i_a(result25[27]), .i_b(~i_divisor[28]), .i_cin(cout26[27]), .i_carry_output(quotient[5]),
		.o_result(result26[28]), .o_cout(cout26[28]));
pu pu26_29 (.i_a(result25[28]), .i_b(~i_divisor[29]), .i_cin(cout26[28]), .i_carry_output(quotient[5]),
		.o_result(result26[29]), .o_cout(cout26[29]));
pu pu26_30 (.i_a(result25[29]), .i_b(~i_divisor[30]), .i_cin(cout26[29]), .i_carry_output(quotient[5]),
		.o_result(result26[30]), .o_cout(cout26[30]));
pu pu26_31 (.i_a(result25[30]), .i_b(~i_divisor[31]), .i_cin(cout26[30]), .i_carry_output(quotient[5]),
		.o_cout(quotient[5]));

// Row 27
pu pu27_0 (.i_a(i_dividend[4]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[4]),
         .o_result(result27[0]), .o_cout(cout27[0]));	
pu pu27_1 (.i_a(result26[0]), .i_b(~i_divisor[1]), .i_cin(cout27[0]), .i_carry_output(quotient[4]),
		.o_result(result27[1]), .o_cout(cout27[1]));
pu pu27_2 (.i_a(result26[1]), .i_b(~i_divisor[2]), .i_cin(cout27[1]), .i_carry_output(quotient[4]),
		.o_result(result27[2]), .o_cout(cout27[2]));
pu pu27_3 (.i_a(result26[2]), .i_b(~i_divisor[3]), .i_cin(cout27[2]), .i_carry_output(quotient[4]),
		.o_result(result27[3]), .o_cout(cout27[3]));
pu pu27_4 (.i_a(result26[3]), .i_b(~i_divisor[4]), .i_cin(cout27[3]), .i_carry_output(quotient[4]),
		.o_result(result27[4]), .o_cout(cout27[4]));
pu pu27_5 (.i_a(result26[4]), .i_b(~i_divisor[5]), .i_cin(cout27[4]), .i_carry_output(quotient[4]),
		.o_result(result27[5]), .o_cout(cout27[5]));
pu pu27_6 (.i_a(result26[5]), .i_b(~i_divisor[6]), .i_cin(cout27[5]), .i_carry_output(quotient[4]),
		.o_result(result27[6]), .o_cout(cout27[6]));
pu pu27_7 (.i_a(result26[6]), .i_b(~i_divisor[7]), .i_cin(cout27[6]), .i_carry_output(quotient[4]),
		.o_result(result27[7]), .o_cout(cout27[7]));
pu pu27_8 (.i_a(result26[7]), .i_b(~i_divisor[8]), .i_cin(cout27[7]), .i_carry_output(quotient[4]),
		.o_result(result27[8]), .o_cout(cout27[8]));
pu pu27_9 (.i_a(result26[8]), .i_b(~i_divisor[9]), .i_cin(cout27[8]), .i_carry_output(quotient[4]),
		.o_result(result27[9]), .o_cout(cout27[9]));
pu pu27_10 (.i_a(result26[9]), .i_b(~i_divisor[10]), .i_cin(cout27[9]), .i_carry_output(quotient[4]),
		.o_result(result27[10]), .o_cout(cout27[10]));
pu pu27_11 (.i_a(result26[10]), .i_b(~i_divisor[11]), .i_cin(cout27[10]), .i_carry_output(quotient[4]),
		.o_result(result27[11]), .o_cout(cout27[11]));
pu pu27_12 (.i_a(result26[11]), .i_b(~i_divisor[12]), .i_cin(cout27[11]), .i_carry_output(quotient[4]),
		.o_result(result27[12]), .o_cout(cout27[12]));
pu pu27_13 (.i_a(result26[12]), .i_b(~i_divisor[13]), .i_cin(cout27[12]), .i_carry_output(quotient[4]),
		.o_result(result27[13]), .o_cout(cout27[13]));
pu pu27_14 (.i_a(result26[13]), .i_b(~i_divisor[14]), .i_cin(cout27[13]), .i_carry_output(quotient[4]),
		.o_result(result27[14]), .o_cout(cout27[14]));
pu pu27_15 (.i_a(result26[14]), .i_b(~i_divisor[15]), .i_cin(cout27[14]), .i_carry_output(quotient[4]),
		.o_result(result27[15]), .o_cout(cout27[15]));
pu pu27_16 (.i_a(result26[15]), .i_b(~i_divisor[16]), .i_cin(cout27[15]), .i_carry_output(quotient[4]),
		.o_result(result27[16]), .o_cout(cout27[16]));
pu pu27_17 (.i_a(result26[16]), .i_b(~i_divisor[17]), .i_cin(cout27[16]), .i_carry_output(quotient[4]),
		.o_result(result27[17]), .o_cout(cout27[17]));
pu pu27_18 (.i_a(result26[17]), .i_b(~i_divisor[18]), .i_cin(cout27[17]), .i_carry_output(quotient[4]),
		.o_result(result27[18]), .o_cout(cout27[18]));
pu pu27_19 (.i_a(result26[18]), .i_b(~i_divisor[19]), .i_cin(cout27[18]), .i_carry_output(quotient[4]),
		.o_result(result27[19]), .o_cout(cout27[19]));
pu pu27_20 (.i_a(result26[19]), .i_b(~i_divisor[20]), .i_cin(cout27[19]), .i_carry_output(quotient[4]),
		.o_result(result27[20]), .o_cout(cout27[20]));
pu pu27_21 (.i_a(result26[20]), .i_b(~i_divisor[21]), .i_cin(cout27[20]), .i_carry_output(quotient[4]),
		.o_result(result27[21]), .o_cout(cout27[21]));
pu pu27_22 (.i_a(result26[21]), .i_b(~i_divisor[22]), .i_cin(cout27[21]), .i_carry_output(quotient[4]),
		.o_result(result27[22]), .o_cout(cout27[22]));
pu pu27_23 (.i_a(result26[22]), .i_b(~i_divisor[23]), .i_cin(cout27[22]), .i_carry_output(quotient[4]),
		.o_result(result27[23]), .o_cout(cout27[23]));
pu pu27_24 (.i_a(result26[23]), .i_b(~i_divisor[24]), .i_cin(cout27[23]), .i_carry_output(quotient[4]),
		.o_result(result27[24]), .o_cout(cout27[24]));
pu pu27_25 (.i_a(result26[24]), .i_b(~i_divisor[25]), .i_cin(cout27[24]), .i_carry_output(quotient[4]),
		.o_result(result27[25]), .o_cout(cout27[25]));
pu pu27_26 (.i_a(result26[25]), .i_b(~i_divisor[26]), .i_cin(cout27[25]), .i_carry_output(quotient[4]),
		.o_result(result27[26]), .o_cout(cout27[26]));
pu pu27_27 (.i_a(result26[26]), .i_b(~i_divisor[27]), .i_cin(cout27[26]), .i_carry_output(quotient[4]),
		.o_result(result27[27]), .o_cout(cout27[27]));
pu pu27_28 (.i_a(result26[27]), .i_b(~i_divisor[28]), .i_cin(cout27[27]), .i_carry_output(quotient[4]),
		.o_result(result27[28]), .o_cout(cout27[28]));
pu pu27_29 (.i_a(result26[28]), .i_b(~i_divisor[29]), .i_cin(cout27[28]), .i_carry_output(quotient[4]),
		.o_result(result27[29]), .o_cout(cout27[29]));
pu pu27_30 (.i_a(result26[29]), .i_b(~i_divisor[30]), .i_cin(cout27[29]), .i_carry_output(quotient[4]),
		.o_result(result27[30]), .o_cout(cout27[30]));
pu pu27_31 (.i_a(result26[30]), .i_b(~i_divisor[31]), .i_cin(cout27[30]), .i_carry_output(quotient[4]),
		.o_cout(quotient[4]));

// Row 28
pu pu28_0 (.i_a(i_dividend[3]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[3]),
         .o_result(result28[0]), .o_cout(cout28[0]));	
pu pu28_1 (.i_a(result27[0]), .i_b(~i_divisor[1]), .i_cin(cout28[0]), .i_carry_output(quotient[3]),
		.o_result(result28[1]), .o_cout(cout28[1]));
pu pu28_2 (.i_a(result27[1]), .i_b(~i_divisor[2]), .i_cin(cout28[1]), .i_carry_output(quotient[3]),
		.o_result(result28[2]), .o_cout(cout28[2]));
pu pu28_3 (.i_a(result27[2]), .i_b(~i_divisor[3]), .i_cin(cout28[2]), .i_carry_output(quotient[3]),
		.o_result(result28[3]), .o_cout(cout28[3]));
pu pu28_4 (.i_a(result27[3]), .i_b(~i_divisor[4]), .i_cin(cout28[3]), .i_carry_output(quotient[3]),
		.o_result(result28[4]), .o_cout(cout28[4]));
pu pu28_5 (.i_a(result27[4]), .i_b(~i_divisor[5]), .i_cin(cout28[4]), .i_carry_output(quotient[3]),
		.o_result(result28[5]), .o_cout(cout28[5]));
pu pu28_6 (.i_a(result27[5]), .i_b(~i_divisor[6]), .i_cin(cout28[5]), .i_carry_output(quotient[3]),
		.o_result(result28[6]), .o_cout(cout28[6]));
pu pu28_7 (.i_a(result27[6]), .i_b(~i_divisor[7]), .i_cin(cout28[6]), .i_carry_output(quotient[3]),
		.o_result(result28[7]), .o_cout(cout28[7]));
pu pu28_8 (.i_a(result27[7]), .i_b(~i_divisor[8]), .i_cin(cout28[7]), .i_carry_output(quotient[3]),
		.o_result(result28[8]), .o_cout(cout28[8]));
pu pu28_9 (.i_a(result27[8]), .i_b(~i_divisor[9]), .i_cin(cout28[8]), .i_carry_output(quotient[3]),
		.o_result(result28[9]), .o_cout(cout28[9]));
pu pu28_10 (.i_a(result27[9]), .i_b(~i_divisor[10]), .i_cin(cout28[9]), .i_carry_output(quotient[3]),
		.o_result(result28[10]), .o_cout(cout28[10]));
pu pu28_11 (.i_a(result27[10]), .i_b(~i_divisor[11]), .i_cin(cout28[10]), .i_carry_output(quotient[3]),
		.o_result(result28[11]), .o_cout(cout28[11]));
pu pu28_12 (.i_a(result27[11]), .i_b(~i_divisor[12]), .i_cin(cout28[11]), .i_carry_output(quotient[3]),
		.o_result(result28[12]), .o_cout(cout28[12]));
pu pu28_13 (.i_a(result27[12]), .i_b(~i_divisor[13]), .i_cin(cout28[12]), .i_carry_output(quotient[3]),
		.o_result(result28[13]), .o_cout(cout28[13]));
pu pu28_14 (.i_a(result27[13]), .i_b(~i_divisor[14]), .i_cin(cout28[13]), .i_carry_output(quotient[3]),
		.o_result(result28[14]), .o_cout(cout28[14]));
pu pu28_15 (.i_a(result27[14]), .i_b(~i_divisor[15]), .i_cin(cout28[14]), .i_carry_output(quotient[3]),
		.o_result(result28[15]), .o_cout(cout28[15]));
pu pu28_16 (.i_a(result27[15]), .i_b(~i_divisor[16]), .i_cin(cout28[15]), .i_carry_output(quotient[3]),
		.o_result(result28[16]), .o_cout(cout28[16]));
pu pu28_17 (.i_a(result27[16]), .i_b(~i_divisor[17]), .i_cin(cout28[16]), .i_carry_output(quotient[3]),
		.o_result(result28[17]), .o_cout(cout28[17]));
pu pu28_18 (.i_a(result27[17]), .i_b(~i_divisor[18]), .i_cin(cout28[17]), .i_carry_output(quotient[3]),
		.o_result(result28[18]), .o_cout(cout28[18]));
pu pu28_19 (.i_a(result27[18]), .i_b(~i_divisor[19]), .i_cin(cout28[18]), .i_carry_output(quotient[3]),
		.o_result(result28[19]), .o_cout(cout28[19]));
pu pu28_20 (.i_a(result27[19]), .i_b(~i_divisor[20]), .i_cin(cout28[19]), .i_carry_output(quotient[3]),
		.o_result(result28[20]), .o_cout(cout28[20]));
pu pu28_21 (.i_a(result27[20]), .i_b(~i_divisor[21]), .i_cin(cout28[20]), .i_carry_output(quotient[3]),
		.o_result(result28[21]), .o_cout(cout28[21]));
pu pu28_22 (.i_a(result27[21]), .i_b(~i_divisor[22]), .i_cin(cout28[21]), .i_carry_output(quotient[3]),
		.o_result(result28[22]), .o_cout(cout28[22]));
pu pu28_23 (.i_a(result27[22]), .i_b(~i_divisor[23]), .i_cin(cout28[22]), .i_carry_output(quotient[3]),
		.o_result(result28[23]), .o_cout(cout28[23]));
pu pu28_24 (.i_a(result27[23]), .i_b(~i_divisor[24]), .i_cin(cout28[23]), .i_carry_output(quotient[3]),
		.o_result(result28[24]), .o_cout(cout28[24]));
pu pu28_25 (.i_a(result27[24]), .i_b(~i_divisor[25]), .i_cin(cout28[24]), .i_carry_output(quotient[3]),
		.o_result(result28[25]), .o_cout(cout28[25]));
pu pu28_26 (.i_a(result27[25]), .i_b(~i_divisor[26]), .i_cin(cout28[25]), .i_carry_output(quotient[3]),
		.o_result(result28[26]), .o_cout(cout28[26]));
pu pu28_27 (.i_a(result27[26]), .i_b(~i_divisor[27]), .i_cin(cout28[26]), .i_carry_output(quotient[3]),
		.o_result(result28[27]), .o_cout(cout28[27]));
pu pu28_28 (.i_a(result27[27]), .i_b(~i_divisor[28]), .i_cin(cout28[27]), .i_carry_output(quotient[3]),
		.o_result(result28[28]), .o_cout(cout28[28]));
pu pu28_29 (.i_a(result27[28]), .i_b(~i_divisor[29]), .i_cin(cout28[28]), .i_carry_output(quotient[3]),
		.o_result(result28[29]), .o_cout(cout28[29]));
pu pu28_30 (.i_a(result27[29]), .i_b(~i_divisor[30]), .i_cin(cout28[29]), .i_carry_output(quotient[3]),
		.o_result(result28[30]), .o_cout(cout28[30]));
pu pu28_31 (.i_a(result27[30]), .i_b(~i_divisor[31]), .i_cin(cout28[30]), .i_carry_output(quotient[3]),
		.o_cout(quotient[3]));

// Row 29
pu pu29_0 (.i_a(i_dividend[2]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[2]),
         .o_result(result29[0]), .o_cout(cout29[0]));	
pu pu29_1 (.i_a(result28[0]), .i_b(~i_divisor[1]), .i_cin(cout29[0]), .i_carry_output(quotient[2]),
		.o_result(result29[1]), .o_cout(cout29[1]));
pu pu29_2 (.i_a(result28[1]), .i_b(~i_divisor[2]), .i_cin(cout29[1]), .i_carry_output(quotient[2]),
		.o_result(result29[2]), .o_cout(cout29[2]));
pu pu29_3 (.i_a(result28[2]), .i_b(~i_divisor[3]), .i_cin(cout29[2]), .i_carry_output(quotient[2]),
		.o_result(result29[3]), .o_cout(cout29[3]));
pu pu29_4 (.i_a(result28[3]), .i_b(~i_divisor[4]), .i_cin(cout29[3]), .i_carry_output(quotient[2]),
		.o_result(result29[4]), .o_cout(cout29[4]));
pu pu29_5 (.i_a(result28[4]), .i_b(~i_divisor[5]), .i_cin(cout29[4]), .i_carry_output(quotient[2]),
		.o_result(result29[5]), .o_cout(cout29[5]));
pu pu29_6 (.i_a(result28[5]), .i_b(~i_divisor[6]), .i_cin(cout29[5]), .i_carry_output(quotient[2]),
		.o_result(result29[6]), .o_cout(cout29[6]));
pu pu29_7 (.i_a(result28[6]), .i_b(~i_divisor[7]), .i_cin(cout29[6]), .i_carry_output(quotient[2]),
		.o_result(result29[7]), .o_cout(cout29[7]));
pu pu29_8 (.i_a(result28[7]), .i_b(~i_divisor[8]), .i_cin(cout29[7]), .i_carry_output(quotient[2]),
		.o_result(result29[8]), .o_cout(cout29[8]));
pu pu29_9 (.i_a(result28[8]), .i_b(~i_divisor[9]), .i_cin(cout29[8]), .i_carry_output(quotient[2]),
		.o_result(result29[9]), .o_cout(cout29[9]));
pu pu29_10 (.i_a(result28[9]), .i_b(~i_divisor[10]), .i_cin(cout29[9]), .i_carry_output(quotient[2]),
		.o_result(result29[10]), .o_cout(cout29[10]));
pu pu29_11 (.i_a(result28[10]), .i_b(~i_divisor[11]), .i_cin(cout29[10]), .i_carry_output(quotient[2]),
		.o_result(result29[11]), .o_cout(cout29[11]));
pu pu29_12 (.i_a(result28[11]), .i_b(~i_divisor[12]), .i_cin(cout29[11]), .i_carry_output(quotient[2]),
		.o_result(result29[12]), .o_cout(cout29[12]));
pu pu29_13 (.i_a(result28[12]), .i_b(~i_divisor[13]), .i_cin(cout29[12]), .i_carry_output(quotient[2]),
		.o_result(result29[13]), .o_cout(cout29[13]));
pu pu29_14 (.i_a(result28[13]), .i_b(~i_divisor[14]), .i_cin(cout29[13]), .i_carry_output(quotient[2]),
		.o_result(result29[14]), .o_cout(cout29[14]));
pu pu29_15 (.i_a(result28[14]), .i_b(~i_divisor[15]), .i_cin(cout29[14]), .i_carry_output(quotient[2]),
		.o_result(result29[15]), .o_cout(cout29[15]));
pu pu29_16 (.i_a(result28[15]), .i_b(~i_divisor[16]), .i_cin(cout29[15]), .i_carry_output(quotient[2]),
		.o_result(result29[16]), .o_cout(cout29[16]));
pu pu29_17 (.i_a(result28[16]), .i_b(~i_divisor[17]), .i_cin(cout29[16]), .i_carry_output(quotient[2]),
		.o_result(result29[17]), .o_cout(cout29[17]));
pu pu29_18 (.i_a(result28[17]), .i_b(~i_divisor[18]), .i_cin(cout29[17]), .i_carry_output(quotient[2]),
		.o_result(result29[18]), .o_cout(cout29[18]));
pu pu29_19 (.i_a(result28[18]), .i_b(~i_divisor[19]), .i_cin(cout29[18]), .i_carry_output(quotient[2]),
		.o_result(result29[19]), .o_cout(cout29[19]));
pu pu29_20 (.i_a(result28[19]), .i_b(~i_divisor[20]), .i_cin(cout29[19]), .i_carry_output(quotient[2]),
		.o_result(result29[20]), .o_cout(cout29[20]));
pu pu29_21 (.i_a(result28[20]), .i_b(~i_divisor[21]), .i_cin(cout29[20]), .i_carry_output(quotient[2]),
		.o_result(result29[21]), .o_cout(cout29[21]));
pu pu29_22 (.i_a(result28[21]), .i_b(~i_divisor[22]), .i_cin(cout29[21]), .i_carry_output(quotient[2]),
		.o_result(result29[22]), .o_cout(cout29[22]));
pu pu29_23 (.i_a(result28[22]), .i_b(~i_divisor[23]), .i_cin(cout29[22]), .i_carry_output(quotient[2]),
		.o_result(result29[23]), .o_cout(cout29[23]));
pu pu29_24 (.i_a(result28[23]), .i_b(~i_divisor[24]), .i_cin(cout29[23]), .i_carry_output(quotient[2]),
		.o_result(result29[24]), .o_cout(cout29[24]));
pu pu29_25 (.i_a(result28[24]), .i_b(~i_divisor[25]), .i_cin(cout29[24]), .i_carry_output(quotient[2]),
		.o_result(result29[25]), .o_cout(cout29[25]));
pu pu29_26 (.i_a(result28[25]), .i_b(~i_divisor[26]), .i_cin(cout29[25]), .i_carry_output(quotient[2]),
		.o_result(result29[26]), .o_cout(cout29[26]));
pu pu29_27 (.i_a(result28[26]), .i_b(~i_divisor[27]), .i_cin(cout29[26]), .i_carry_output(quotient[2]),
		.o_result(result29[27]), .o_cout(cout29[27]));
pu pu29_28 (.i_a(result28[27]), .i_b(~i_divisor[28]), .i_cin(cout29[27]), .i_carry_output(quotient[2]),
		.o_result(result29[28]), .o_cout(cout29[28]));
pu pu29_29 (.i_a(result28[28]), .i_b(~i_divisor[29]), .i_cin(cout29[28]), .i_carry_output(quotient[2]),
		.o_result(result29[29]), .o_cout(cout29[29]));
pu pu29_30 (.i_a(result28[29]), .i_b(~i_divisor[30]), .i_cin(cout29[29]), .i_carry_output(quotient[2]),
		.o_result(result29[30]), .o_cout(cout29[30]));
pu pu29_31 (.i_a(result28[30]), .i_b(~i_divisor[31]), .i_cin(cout29[30]), .i_carry_output(quotient[2]),
		.o_cout(quotient[2]));

// Row 30
pu pu30_0 (.i_a(i_dividend[1]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[1]),
         .o_result(result30[0]), .o_cout(cout30[0]));	
pu pu30_1 (.i_a(result29[0]), .i_b(~i_divisor[1]), .i_cin(cout30[0]), .i_carry_output(quotient[1]),
		.o_result(result30[1]), .o_cout(cout30[1]));
pu pu30_2 (.i_a(result29[1]), .i_b(~i_divisor[2]), .i_cin(cout30[1]), .i_carry_output(quotient[1]),
		.o_result(result30[2]), .o_cout(cout30[2]));
pu pu30_3 (.i_a(result29[2]), .i_b(~i_divisor[3]), .i_cin(cout30[2]), .i_carry_output(quotient[1]),
		.o_result(result30[3]), .o_cout(cout30[3]));
pu pu30_4 (.i_a(result29[3]), .i_b(~i_divisor[4]), .i_cin(cout30[3]), .i_carry_output(quotient[1]),
		.o_result(result30[4]), .o_cout(cout30[4]));
pu pu30_5 (.i_a(result29[4]), .i_b(~i_divisor[5]), .i_cin(cout30[4]), .i_carry_output(quotient[1]),
		.o_result(result30[5]), .o_cout(cout30[5]));
pu pu30_6 (.i_a(result29[5]), .i_b(~i_divisor[6]), .i_cin(cout30[5]), .i_carry_output(quotient[1]),
		.o_result(result30[6]), .o_cout(cout30[6]));
pu pu30_7 (.i_a(result29[6]), .i_b(~i_divisor[7]), .i_cin(cout30[6]), .i_carry_output(quotient[1]),
		.o_result(result30[7]), .o_cout(cout30[7]));
pu pu30_8 (.i_a(result29[7]), .i_b(~i_divisor[8]), .i_cin(cout30[7]), .i_carry_output(quotient[1]),
		.o_result(result30[8]), .o_cout(cout30[8]));
pu pu30_9 (.i_a(result29[8]), .i_b(~i_divisor[9]), .i_cin(cout30[8]), .i_carry_output(quotient[1]),
		.o_result(result30[9]), .o_cout(cout30[9]));
pu pu30_10 (.i_a(result29[9]), .i_b(~i_divisor[10]), .i_cin(cout30[9]), .i_carry_output(quotient[1]),
		.o_result(result30[10]), .o_cout(cout30[10]));
pu pu30_11 (.i_a(result29[10]), .i_b(~i_divisor[11]), .i_cin(cout30[10]), .i_carry_output(quotient[1]),
		.o_result(result30[11]), .o_cout(cout30[11]));
pu pu30_12 (.i_a(result29[11]), .i_b(~i_divisor[12]), .i_cin(cout30[11]), .i_carry_output(quotient[1]),
		.o_result(result30[12]), .o_cout(cout30[12]));
pu pu30_13 (.i_a(result29[12]), .i_b(~i_divisor[13]), .i_cin(cout30[12]), .i_carry_output(quotient[1]),
		.o_result(result30[13]), .o_cout(cout30[13]));
pu pu30_14 (.i_a(result29[13]), .i_b(~i_divisor[14]), .i_cin(cout30[13]), .i_carry_output(quotient[1]),
		.o_result(result30[14]), .o_cout(cout30[14]));
pu pu30_15 (.i_a(result29[14]), .i_b(~i_divisor[15]), .i_cin(cout30[14]), .i_carry_output(quotient[1]),
		.o_result(result30[15]), .o_cout(cout30[15]));
pu pu30_16 (.i_a(result29[15]), .i_b(~i_divisor[16]), .i_cin(cout30[15]), .i_carry_output(quotient[1]),
		.o_result(result30[16]), .o_cout(cout30[16]));
pu pu30_17 (.i_a(result29[16]), .i_b(~i_divisor[17]), .i_cin(cout30[16]), .i_carry_output(quotient[1]),
		.o_result(result30[17]), .o_cout(cout30[17]));
pu pu30_18 (.i_a(result29[17]), .i_b(~i_divisor[18]), .i_cin(cout30[17]), .i_carry_output(quotient[1]),
		.o_result(result30[18]), .o_cout(cout30[18]));
pu pu30_19 (.i_a(result29[18]), .i_b(~i_divisor[19]), .i_cin(cout30[18]), .i_carry_output(quotient[1]),
		.o_result(result30[19]), .o_cout(cout30[19]));
pu pu30_20 (.i_a(result29[19]), .i_b(~i_divisor[20]), .i_cin(cout30[19]), .i_carry_output(quotient[1]),
		.o_result(result30[20]), .o_cout(cout30[20]));
pu pu30_21 (.i_a(result29[20]), .i_b(~i_divisor[21]), .i_cin(cout30[20]), .i_carry_output(quotient[1]),
		.o_result(result30[21]), .o_cout(cout30[21]));
pu pu30_22 (.i_a(result29[21]), .i_b(~i_divisor[22]), .i_cin(cout30[21]), .i_carry_output(quotient[1]),
		.o_result(result30[22]), .o_cout(cout30[22]));
pu pu30_23 (.i_a(result29[22]), .i_b(~i_divisor[23]), .i_cin(cout30[22]), .i_carry_output(quotient[1]),
		.o_result(result30[23]), .o_cout(cout30[23]));
pu pu30_24 (.i_a(result29[23]), .i_b(~i_divisor[24]), .i_cin(cout30[23]), .i_carry_output(quotient[1]),
		.o_result(result30[24]), .o_cout(cout30[24]));
pu pu30_25 (.i_a(result29[24]), .i_b(~i_divisor[25]), .i_cin(cout30[24]), .i_carry_output(quotient[1]),
		.o_result(result30[25]), .o_cout(cout30[25]));
pu pu30_26 (.i_a(result29[25]), .i_b(~i_divisor[26]), .i_cin(cout30[25]), .i_carry_output(quotient[1]),
		.o_result(result30[26]), .o_cout(cout30[26]));
pu pu30_27 (.i_a(result29[26]), .i_b(~i_divisor[27]), .i_cin(cout30[26]), .i_carry_output(quotient[1]),
		.o_result(result30[27]), .o_cout(cout30[27]));
pu pu30_28 (.i_a(result29[27]), .i_b(~i_divisor[28]), .i_cin(cout30[27]), .i_carry_output(quotient[1]),
		.o_result(result30[28]), .o_cout(cout30[28]));
pu pu30_29 (.i_a(result29[28]), .i_b(~i_divisor[29]), .i_cin(cout30[28]), .i_carry_output(quotient[1]),
		.o_result(result30[29]), .o_cout(cout30[29]));
pu pu30_30 (.i_a(result29[29]), .i_b(~i_divisor[30]), .i_cin(cout30[29]), .i_carry_output(quotient[1]),
		.o_result(result30[30]), .o_cout(cout30[30]));
pu pu30_31 (.i_a(result29[30]), .i_b(~i_divisor[31]), .i_cin(cout30[30]), .i_carry_output(quotient[1]),
		.o_cout(quotient[1]));

// Row 31
pu pu31_0 (.i_a(i_dividend[0]), .i_b(~i_divisor[0]), .i_cin(1), .i_carry_output(quotient[0]),
         .o_result(result31[0]), .o_cout(cout31[0]));	
pu pu31_1 (.i_a(result30[0]), .i_b(~i_divisor[1]), .i_cin(cout31[0]), .i_carry_output(quotient[0]),
		.o_result(result31[1]), .o_cout(cout31[1]));
pu pu31_2 (.i_a(result30[1]), .i_b(~i_divisor[2]), .i_cin(cout31[1]), .i_carry_output(quotient[0]),
		.o_result(result31[2]), .o_cout(cout31[2]));
pu pu31_3 (.i_a(result30[2]), .i_b(~i_divisor[3]), .i_cin(cout31[2]), .i_carry_output(quotient[0]),
		.o_result(result31[3]), .o_cout(cout31[3]));
pu pu31_4 (.i_a(result30[3]), .i_b(~i_divisor[4]), .i_cin(cout31[3]), .i_carry_output(quotient[0]),
		.o_result(result31[4]), .o_cout(cout31[4]));
pu pu31_5 (.i_a(result30[4]), .i_b(~i_divisor[5]), .i_cin(cout31[4]), .i_carry_output(quotient[0]),
		.o_result(result31[5]), .o_cout(cout31[5]));
pu pu31_6 (.i_a(result30[5]), .i_b(~i_divisor[6]), .i_cin(cout31[5]), .i_carry_output(quotient[0]),
		.o_result(result31[6]), .o_cout(cout31[6]));
pu pu31_7 (.i_a(result30[6]), .i_b(~i_divisor[7]), .i_cin(cout31[6]), .i_carry_output(quotient[0]),
		.o_result(result31[7]), .o_cout(cout31[7]));
pu pu31_8 (.i_a(result30[7]), .i_b(~i_divisor[8]), .i_cin(cout31[7]), .i_carry_output(quotient[0]),
		.o_result(result31[8]), .o_cout(cout31[8]));
pu pu31_9 (.i_a(result30[8]), .i_b(~i_divisor[9]), .i_cin(cout31[8]), .i_carry_output(quotient[0]),
		.o_result(result31[9]), .o_cout(cout31[9]));
pu pu31_10 (.i_a(result30[9]), .i_b(~i_divisor[10]), .i_cin(cout31[9]), .i_carry_output(quotient[0]),
		.o_result(result31[10]), .o_cout(cout31[10]));
pu pu31_11 (.i_a(result30[10]), .i_b(~i_divisor[11]), .i_cin(cout31[10]), .i_carry_output(quotient[0]),
		.o_result(result31[11]), .o_cout(cout31[11]));
pu pu31_12 (.i_a(result30[11]), .i_b(~i_divisor[12]), .i_cin(cout31[11]), .i_carry_output(quotient[0]),
		.o_result(result31[12]), .o_cout(cout31[12]));
pu pu31_13 (.i_a(result30[12]), .i_b(~i_divisor[13]), .i_cin(cout31[12]), .i_carry_output(quotient[0]),
		.o_result(result31[13]), .o_cout(cout31[13]));
pu pu31_14 (.i_a(result30[13]), .i_b(~i_divisor[14]), .i_cin(cout31[13]), .i_carry_output(quotient[0]),
		.o_result(result31[14]), .o_cout(cout31[14]));
pu pu31_15 (.i_a(result30[14]), .i_b(~i_divisor[15]), .i_cin(cout31[14]), .i_carry_output(quotient[0]),
		.o_result(result31[15]), .o_cout(cout31[15]));
pu pu31_16 (.i_a(result30[15]), .i_b(~i_divisor[16]), .i_cin(cout31[15]), .i_carry_output(quotient[0]),
		.o_result(result31[16]), .o_cout(cout31[16]));
pu pu31_17 (.i_a(result30[16]), .i_b(~i_divisor[17]), .i_cin(cout31[16]), .i_carry_output(quotient[0]),
		.o_result(result31[17]), .o_cout(cout31[17]));
pu pu31_18 (.i_a(result30[17]), .i_b(~i_divisor[18]), .i_cin(cout31[17]), .i_carry_output(quotient[0]),
		.o_result(result31[18]), .o_cout(cout31[18]));
pu pu31_19 (.i_a(result30[18]), .i_b(~i_divisor[19]), .i_cin(cout31[18]), .i_carry_output(quotient[0]),
		.o_result(result31[19]), .o_cout(cout31[19]));
pu pu31_20 (.i_a(result30[19]), .i_b(~i_divisor[20]), .i_cin(cout31[19]), .i_carry_output(quotient[0]),
		.o_result(result31[20]), .o_cout(cout31[20]));
pu pu31_21 (.i_a(result30[20]), .i_b(~i_divisor[21]), .i_cin(cout31[20]), .i_carry_output(quotient[0]),
		.o_result(result31[21]), .o_cout(cout31[21]));
pu pu31_22 (.i_a(result30[21]), .i_b(~i_divisor[22]), .i_cin(cout31[21]), .i_carry_output(quotient[0]),
		.o_result(result31[22]), .o_cout(cout31[22]));
pu pu31_23 (.i_a(result30[22]), .i_b(~i_divisor[23]), .i_cin(cout31[22]), .i_carry_output(quotient[0]),
		.o_result(result31[23]), .o_cout(cout31[23]));
pu pu31_24 (.i_a(result30[23]), .i_b(~i_divisor[24]), .i_cin(cout31[23]), .i_carry_output(quotient[0]),
		.o_result(result31[24]), .o_cout(cout31[24]));
pu pu31_25 (.i_a(result30[24]), .i_b(~i_divisor[25]), .i_cin(cout31[24]), .i_carry_output(quotient[0]),
		.o_result(result31[25]), .o_cout(cout31[25]));
pu pu31_26 (.i_a(result30[25]), .i_b(~i_divisor[26]), .i_cin(cout31[25]), .i_carry_output(quotient[0]),
		.o_result(result31[26]), .o_cout(cout31[26]));
pu pu31_27 (.i_a(result30[26]), .i_b(~i_divisor[27]), .i_cin(cout31[26]), .i_carry_output(quotient[0]),
		.o_result(result31[27]), .o_cout(cout31[27]));
pu pu31_28 (.i_a(result30[27]), .i_b(~i_divisor[28]), .i_cin(cout31[27]), .i_carry_output(quotient[0]),
		.o_result(result31[28]), .o_cout(cout31[28]));
pu pu31_29 (.i_a(result30[28]), .i_b(~i_divisor[29]), .i_cin(cout31[28]), .i_carry_output(quotient[0]),
		.o_result(result31[29]), .o_cout(cout31[29]));
pu pu31_30 (.i_a(result30[29]), .i_b(~i_divisor[30]), .i_cin(cout31[29]), .i_carry_output(quotient[0]),
		.o_result(result31[30]), .o_cout(cout31[30]));
pu pu31_31 (.i_a(result30[30]), .i_b(~i_divisor[31]), .i_cin(cout31[30]), .i_carry_output(quotient[0]),
		.o_result(result31[31]), .o_cout(quotient[0]));

always @(*) begin
	if (i_divisor == 32'b0) begin
		o_quotient = 32'hFFFF_FFFF;
		o_remainder = i_dividend;
	end else begin
		o_remainder = result31;
		o_quotient = quotient;
	end
end

endmodule

module pu (
	input logic i_a, i_b, i_cin, i_carry_output,
	output logic o_result, o_cout
);

logic sum;

fullAdder fa1 (.a(i_a), .b(i_b), .cin(i_cin), .cout(o_cout), .sum(sum));

always @(*) begin
	if (i_carry_output) 
		o_result = sum;
	else
		o_result = i_a;
end

endmodule
