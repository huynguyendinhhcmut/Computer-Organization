/*
==================================================================================================
		 ___                      ____            
		|_ _|_ __ ___  _ __ ___  / ___| ___ _ __  
		 | || '_ ` _ \| '_ ` _ \| |  _ / _ \ '_ \ 
		 | || | | | | | | | | | | |_| |  __/ | | |
		|___|_| |_| |_|_| |_| |_|\____|\___|_| |_|
                                                        
==================================================================================================
*/
module ImmGen 
(
	input	[24:0]	instr,			// Range contaim Immediate [31:7]
	input [2:0]		imm_sel,			// Select which range contain Immediate			// Select Size and Signed or not
	output[31:0]	ImmExt			// Output of full Immediate
);

/*

	|--------------------|-----------|-----------|-----------|-----------|-----------------------------------------------------------------|
	|	 	Description		| imm_sel2	| imm_sel1	|	imm_sel0	|	  Type 	|										Imm Ext										|
	|--------------------|-----------|-----------|-----------|-----------|-----------------------------------------------------------------|
	|		12-bit signed	|		0		|		0		|		0		|		I		|						 {{20{Instr[31]}}, Instr[31:20]}						|
	|--------------------|-----------|-----------|-----------|-----------|-----------------------------------------------------------------|
	|		12-bit signed	|		0		|		0		|		1		|		S		|			{{20{Instr[31]}}, Instr[31:25], Instr[11:7]}					|
	|--------------------|-----------|-----------|-----------|-----------|-----------------------------------------------------------------|
	|		12-bit signed	|		0		|		1		|		0		|		B		|	{{20{Instr[31]}}, Instr[7], Instr[30:25], Instr[11:8], 1’b0}	|
	|--------------------|-----------|-----------|-----------|-----------|-----------------------------------------------------------------|
	|		21-bit signed 	|		0		|		1		|		1		|		J		|  {{12{Instr[31]}}, Instr[19:12], Instr[20], Instr[30:21], 1’b0} |
	|--------------------|-----------|-----------|-----------|-----------|-----------------------------------------------------------------|
	|		20-bit signed	|		1		|		0		|		0		|		U		|							  {Instr[31:12], 12'b0}								|
	|--------------------|-----------|-----------|-----------|-----------|-----------------------------------------------------------------|
	
*/

always @(*) begin
    case (imm_sel)
		3'b000: ImmExt = {{20{instr[24]}}, instr[24:13]};												// I Type
		3'b001: ImmExt = {{20{instr[24]}}, instr[24:18], instr[4:0]};								// S Type
		3'b010: ImmExt = {{20{instr[24]}}, instr[0], instr[23:18], instr[4:1], 1'b0};			// B Type
		3'b011: ImmExt = {{12{instr[24]}}, instr[12:5], instr[13], instr[23:14], 1'b0};		// J Type
		3'b100: ImmExt = {instr[24:5], 12'b0};																// U Type
		default: ImmExt = 32'b0;
	endcase
end



endmodule 



