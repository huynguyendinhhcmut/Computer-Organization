module ram_tag_valid (
    input logic  i_clk,
    input logic  i_btb_wren,
    input logic  [9:0]  i_addr,
    input logic  [31:0] i_data,
    
	output logic [31:0] o_data
);

reg [31:0] ram [0:1023];

initial begin
        $readmemh("/home/yellow/ctmt_cttt_4/pipelined_fowarding_g_share/02_test/bht_init_file.hex", ram);
end

always_ff @(posedge i_clk) begin
	if (i_btb_wren) begin
		ram[i_addr] <= i_data;
	end
end

always_ff @(negedge i_clk) begin
	o_data <= ram[i_addr];
end

endmodule

