module instrmem (
    input  logic [31:0] i_pc,
    output logic [31:0] o_instr
);

logic [3:0][7:0] memory [0:1999];  
logic [7:0] temp_mem [0:7999];   
	
initial begin
   $readmemh("program.txt", temp_mem);

   memory[0][0] = temp_mem[0];
   memory[0][1] = temp_mem[1];
   memory[0][2] = temp_mem[2];
   memory[0][3] = temp_mem[3];

   memory[1][0] = temp_mem[4];
   memory[1][1] = temp_mem[5];
   memory[1][2] = temp_mem[6];
   memory[1][3] = temp_mem[7];

   memory[2][0] = temp_mem[8];
   memory[2][1] = temp_mem[9];
   memory[2][2] = temp_mem[10];
   memory[2][3] = temp_mem[11];

   memory[3][0] = temp_mem[12];
   memory[3][1] = temp_mem[13];
   memory[3][2] = temp_mem[14];
   memory[3][3] = temp_mem[15];

   memory[4][0] = temp_mem[16];
   memory[4][1] = temp_mem[17];
   memory[4][2] = temp_mem[18];
   memory[4][3] = temp_mem[19];

   memory[5][0] = temp_mem[20];
   memory[5][1] = temp_mem[21];
   memory[5][2] = temp_mem[22];
   memory[5][3] = temp_mem[23];

   memory[6][0] = temp_mem[24];
   memory[6][1] = temp_mem[25];
   memory[6][2] = temp_mem[26];
   memory[6][3] = temp_mem[27];

   memory[7][0] = temp_mem[28];
   memory[7][1] = temp_mem[29];
   memory[7][2] = temp_mem[30];
   memory[7][3] = temp_mem[31];

   memory[8][0] = temp_mem[32];
   memory[8][1] = temp_mem[33];
   memory[8][2] = temp_mem[34];
   memory[8][3] = temp_mem[35];

   memory[9][0] = temp_mem[36];
   memory[9][1] = temp_mem[37];
   memory[9][2] = temp_mem[38];
   memory[9][3] = temp_mem[39];

   memory[10][0] = temp_mem[40];
   memory[10][1] = temp_mem[41];
   memory[10][2] = temp_mem[42];
   memory[10][3] = temp_mem[43];

   memory[11][0] = temp_mem[44];
   memory[11][1] = temp_mem[45];
   memory[11][2] = temp_mem[46];
   memory[11][3] = temp_mem[47];

   memory[12][0] = temp_mem[48];
   memory[12][1] = temp_mem[49];
   memory[12][2] = temp_mem[50];
   memory[12][3] = temp_mem[51];

   memory[13][0] = temp_mem[52];
   memory[13][1] = temp_mem[53];
   memory[13][2] = temp_mem[54];
   memory[13][3] = temp_mem[55];

   memory[14][0] = temp_mem[56];
   memory[14][1] = temp_mem[57];
   memory[14][2] = temp_mem[58];
   memory[14][3] = temp_mem[59];

   memory[15][0] = temp_mem[60];
   memory[15][1] = temp_mem[61];
   memory[15][2] = temp_mem[62];
   memory[15][3] = temp_mem[63];

   memory[16][0] = temp_mem[64];
   memory[16][1] = temp_mem[65];
   memory[16][2] = temp_mem[66];
   memory[16][3] = temp_mem[67];

   memory[17][0] = temp_mem[68];
   memory[17][1] = temp_mem[69];
   memory[17][2] = temp_mem[70];
   memory[17][3] = temp_mem[71];

   memory[18][0] = temp_mem[72];
   memory[18][1] = temp_mem[73];
   memory[18][2] = temp_mem[74];
   memory[18][3] = temp_mem[75];

   memory[19][0] = temp_mem[76];
   memory[19][1] = temp_mem[77];
   memory[19][2] = temp_mem[78];
   memory[19][3] = temp_mem[79];

   memory[20][0] = temp_mem[80];
   memory[20][1] = temp_mem[81];
   memory[20][2] = temp_mem[82];
   memory[20][3] = temp_mem[83];

   memory[21][0] = temp_mem[84];
   memory[21][1] = temp_mem[85];
   memory[21][2] = temp_mem[86];
   memory[21][3] = temp_mem[87];

   memory[22][0] = temp_mem[88];
   memory[22][1] = temp_mem[89];
   memory[22][2] = temp_mem[90];
   memory[22][3] = temp_mem[91];

   memory[23][0] = temp_mem[92];
   memory[23][1] = temp_mem[93];
   memory[23][2] = temp_mem[94];
   memory[23][3] = temp_mem[95];

   memory[24][0] = temp_mem[96];
   memory[24][1] = temp_mem[97];
   memory[24][2] = temp_mem[98];
   memory[24][3] = temp_mem[99];

   memory[25][0] = temp_mem[100];
   memory[25][1] = temp_mem[101];
   memory[25][2] = temp_mem[102];
   memory[25][3] = temp_mem[103];

   memory[26][0] = temp_mem[104];
   memory[26][1] = temp_mem[105];
   memory[26][2] = temp_mem[106];
   memory[26][3] = temp_mem[107];

   memory[27][0] = temp_mem[108];
   memory[27][1] = temp_mem[109];
   memory[27][2] = temp_mem[110];
   memory[27][3] = temp_mem[111];

   memory[28][0] = temp_mem[112];
   memory[28][1] = temp_mem[113];
   memory[28][2] = temp_mem[114];
   memory[28][3] = temp_mem[115];

   memory[29][0] = temp_mem[116];
   memory[29][1] = temp_mem[117];
   memory[29][2] = temp_mem[118];
   memory[29][3] = temp_mem[119];

   memory[30][0] = temp_mem[120];
   memory[30][1] = temp_mem[121];
   memory[30][2] = temp_mem[122];
   memory[30][3] = temp_mem[123];

   memory[31][0] = temp_mem[124];
   memory[31][1] = temp_mem[125];
   memory[31][2] = temp_mem[126];
   memory[31][3] = temp_mem[127];

   memory[32][0] = temp_mem[128];
   memory[32][1] = temp_mem[129];
   memory[32][2] = temp_mem[130];
   memory[32][3] = temp_mem[131];

   memory[33][0] = temp_mem[132];
   memory[33][1] = temp_mem[133];
   memory[33][2] = temp_mem[134];
   memory[33][3] = temp_mem[135];

   memory[34][0] = temp_mem[136];
   memory[34][1] = temp_mem[137];
   memory[34][2] = temp_mem[138];
   memory[34][3] = temp_mem[139];

   memory[35][0] = temp_mem[140];
   memory[35][1] = temp_mem[141];
   memory[35][2] = temp_mem[142];
   memory[35][3] = temp_mem[143];

   memory[36][0] = temp_mem[144];
   memory[36][1] = temp_mem[145];
   memory[36][2] = temp_mem[146];
   memory[36][3] = temp_mem[147];

   memory[37][0] = temp_mem[148];
   memory[37][1] = temp_mem[149];
   memory[37][2] = temp_mem[150];
   memory[37][3] = temp_mem[151];

   memory[38][0] = temp_mem[152];
   memory[38][1] = temp_mem[153];
   memory[38][2] = temp_mem[154];
   memory[38][3] = temp_mem[155];

   memory[39][0] = temp_mem[156];
   memory[39][1] = temp_mem[157];
   memory[39][2] = temp_mem[158];
   memory[39][3] = temp_mem[159];

   memory[40][0] = temp_mem[160];
   memory[40][1] = temp_mem[161];
   memory[40][2] = temp_mem[162];
   memory[40][3] = temp_mem[163];

   memory[41][0] = temp_mem[164];
   memory[41][1] = temp_mem[165];
   memory[41][2] = temp_mem[166];
   memory[41][3] = temp_mem[167];

   memory[42][0] = temp_mem[168];
   memory[42][1] = temp_mem[169];
   memory[42][2] = temp_mem[170];
   memory[42][3] = temp_mem[171];

   memory[43][0] = temp_mem[172];
   memory[43][1] = temp_mem[173];
   memory[43][2] = temp_mem[174];
   memory[43][3] = temp_mem[175];

   memory[44][0] = temp_mem[176];
   memory[44][1] = temp_mem[177];
   memory[44][2] = temp_mem[178];
   memory[44][3] = temp_mem[179];

   memory[45][0] = temp_mem[180];
   memory[45][1] = temp_mem[181];
   memory[45][2] = temp_mem[182];
   memory[45][3] = temp_mem[183];

   memory[46][0] = temp_mem[184];
   memory[46][1] = temp_mem[185];
   memory[46][2] = temp_mem[186];
   memory[46][3] = temp_mem[187];

   memory[47][0] = temp_mem[188];
   memory[47][1] = temp_mem[189];
   memory[47][2] = temp_mem[190];
   memory[47][3] = temp_mem[191];

   memory[48][0] = temp_mem[192];
   memory[48][1] = temp_mem[193];
   memory[48][2] = temp_mem[194];
   memory[48][3] = temp_mem[195];

   memory[49][0] = temp_mem[196];
   memory[49][1] = temp_mem[197];
   memory[49][2] = temp_mem[198];
   memory[49][3] = temp_mem[199];

   memory[50][0] = temp_mem[200];
   memory[50][1] = temp_mem[201];
   memory[50][2] = temp_mem[202];
   memory[50][3] = temp_mem[203];

   memory[51][0] = temp_mem[204];
   memory[51][1] = temp_mem[205];
   memory[51][2] = temp_mem[206];
   memory[51][3] = temp_mem[207];

   memory[52][0] = temp_mem[208];
   memory[52][1] = temp_mem[209];
   memory[52][2] = temp_mem[210];
   memory[52][3] = temp_mem[211];

   memory[53][0] = temp_mem[212];
   memory[53][1] = temp_mem[213];
   memory[53][2] = temp_mem[214];
   memory[53][3] = temp_mem[215];

   memory[54][0] = temp_mem[216];
   memory[54][1] = temp_mem[217];
   memory[54][2] = temp_mem[218];
   memory[54][3] = temp_mem[219];

   memory[55][0] = temp_mem[220];
   memory[55][1] = temp_mem[221];
   memory[55][2] = temp_mem[222];
   memory[55][3] = temp_mem[223];

   memory[56][0] = temp_mem[224];
   memory[56][1] = temp_mem[225];
   memory[56][2] = temp_mem[226];
   memory[56][3] = temp_mem[227];

   memory[57][0] = temp_mem[228];
   memory[57][1] = temp_mem[229];
   memory[57][2] = temp_mem[230];
   memory[57][3] = temp_mem[231];

   memory[58][0] = temp_mem[232];
   memory[58][1] = temp_mem[233];
   memory[58][2] = temp_mem[234];
   memory[58][3] = temp_mem[235];

   memory[59][0] = temp_mem[236];
   memory[59][1] = temp_mem[237];
   memory[59][2] = temp_mem[238];
   memory[59][3] = temp_mem[239];

   memory[60][0] = temp_mem[240];
   memory[60][1] = temp_mem[241];
   memory[60][2] = temp_mem[242];
   memory[60][3] = temp_mem[243];

   memory[61][0] = temp_mem[244];
   memory[61][1] = temp_mem[245];
   memory[61][2] = temp_mem[246];
   memory[61][3] = temp_mem[247];

   memory[62][0] = temp_mem[248];
   memory[62][1] = temp_mem[249];
   memory[62][2] = temp_mem[250];
   memory[62][3] = temp_mem[251];

   memory[63][0] = temp_mem[252];
   memory[63][1] = temp_mem[253];
   memory[63][2] = temp_mem[254];
   memory[63][3] = temp_mem[255];

   memory[64][0] = temp_mem[256];
   memory[64][1] = temp_mem[257];
   memory[64][2] = temp_mem[258];
   memory[64][3] = temp_mem[259];

   memory[65][0] = temp_mem[260];
   memory[65][1] = temp_mem[261];
   memory[65][2] = temp_mem[262];
   memory[65][3] = temp_mem[263];

   memory[66][0] = temp_mem[264];
   memory[66][1] = temp_mem[265];
   memory[66][2] = temp_mem[266];
   memory[66][3] = temp_mem[267];

   memory[67][0] = temp_mem[268];
   memory[67][1] = temp_mem[269];
   memory[67][2] = temp_mem[270];
   memory[67][3] = temp_mem[271];

   memory[68][0] = temp_mem[272];
   memory[68][1] = temp_mem[273];
   memory[68][2] = temp_mem[274];
   memory[68][3] = temp_mem[275];

   memory[69][0] = temp_mem[276];
   memory[69][1] = temp_mem[277];
   memory[69][2] = temp_mem[278];
   memory[69][3] = temp_mem[279];

   memory[70][0] = temp_mem[280];
   memory[70][1] = temp_mem[281];
   memory[70][2] = temp_mem[282];
   memory[70][3] = temp_mem[283];

   memory[71][0] = temp_mem[284];
   memory[71][1] = temp_mem[285];
   memory[71][2] = temp_mem[286];
   memory[71][3] = temp_mem[287];

   memory[72][0] = temp_mem[288];
   memory[72][1] = temp_mem[289];
   memory[72][2] = temp_mem[290];
   memory[72][3] = temp_mem[291];

   memory[73][0] = temp_mem[292];
   memory[73][1] = temp_mem[293];
   memory[73][2] = temp_mem[294];
   memory[73][3] = temp_mem[295];

   memory[74][0] = temp_mem[296];
   memory[74][1] = temp_mem[297];
   memory[74][2] = temp_mem[298];
   memory[74][3] = temp_mem[299];

   memory[75][0] = temp_mem[300];
   memory[75][1] = temp_mem[301];
   memory[75][2] = temp_mem[302];
   memory[75][3] = temp_mem[303];

   memory[76][0] = temp_mem[304];
   memory[76][1] = temp_mem[305];
   memory[76][2] = temp_mem[306];
   memory[76][3] = temp_mem[307];

   memory[77][0] = temp_mem[308];
   memory[77][1] = temp_mem[309];
   memory[77][2] = temp_mem[310];
   memory[77][3] = temp_mem[311];

   memory[78][0] = temp_mem[312];
   memory[78][1] = temp_mem[313];
   memory[78][2] = temp_mem[314];
   memory[78][3] = temp_mem[315];

   memory[79][0] = temp_mem[316];
   memory[79][1] = temp_mem[317];
   memory[79][2] = temp_mem[318];
   memory[79][3] = temp_mem[319];

   memory[80][0] = temp_mem[320];
   memory[80][1] = temp_mem[321];
   memory[80][2] = temp_mem[322];
   memory[80][3] = temp_mem[323];

   memory[81][0] = temp_mem[324];
   memory[81][1] = temp_mem[325];
   memory[81][2] = temp_mem[326];
   memory[81][3] = temp_mem[327];

   memory[82][0] = temp_mem[328];
   memory[82][1] = temp_mem[329];
   memory[82][2] = temp_mem[330];
   memory[82][3] = temp_mem[331];

   memory[83][0] = temp_mem[332];
   memory[83][1] = temp_mem[333];
   memory[83][2] = temp_mem[334];
   memory[83][3] = temp_mem[335];

   memory[84][0] = temp_mem[336];
   memory[84][1] = temp_mem[337];
   memory[84][2] = temp_mem[338];
   memory[84][3] = temp_mem[339];

   memory[85][0] = temp_mem[340];
   memory[85][1] = temp_mem[341];
   memory[85][2] = temp_mem[342];
   memory[85][3] = temp_mem[343];

   memory[86][0] = temp_mem[344];
   memory[86][1] = temp_mem[345];
   memory[86][2] = temp_mem[346];
   memory[86][3] = temp_mem[347];

   memory[87][0] = temp_mem[348];
   memory[87][1] = temp_mem[349];
   memory[87][2] = temp_mem[350];
   memory[87][3] = temp_mem[351];

   memory[88][0] = temp_mem[352];
   memory[88][1] = temp_mem[353];
   memory[88][2] = temp_mem[354];
   memory[88][3] = temp_mem[355];

   memory[89][0] = temp_mem[356];
   memory[89][1] = temp_mem[357];
   memory[89][2] = temp_mem[358];
   memory[89][3] = temp_mem[359];

   memory[90][0] = temp_mem[360];
   memory[90][1] = temp_mem[361];
   memory[90][2] = temp_mem[362];
   memory[90][3] = temp_mem[363];

   memory[91][0] = temp_mem[364];
   memory[91][1] = temp_mem[365];
   memory[91][2] = temp_mem[366];
   memory[91][3] = temp_mem[367];

   memory[92][0] = temp_mem[368];
   memory[92][1] = temp_mem[369];
   memory[92][2] = temp_mem[370];
   memory[92][3] = temp_mem[371];

   memory[93][0] = temp_mem[372];
   memory[93][1] = temp_mem[373];
   memory[93][2] = temp_mem[374];
   memory[93][3] = temp_mem[375];

   memory[94][0] = temp_mem[376];
   memory[94][1] = temp_mem[377];
   memory[94][2] = temp_mem[378];
   memory[94][3] = temp_mem[379];

   memory[95][0] = temp_mem[380];
   memory[95][1] = temp_mem[381];
   memory[95][2] = temp_mem[382];
   memory[95][3] = temp_mem[383];

   memory[96][0] = temp_mem[384];
   memory[96][1] = temp_mem[385];
   memory[96][2] = temp_mem[386];
   memory[96][3] = temp_mem[387];

   memory[97][0] = temp_mem[388];
   memory[97][1] = temp_mem[389];
   memory[97][2] = temp_mem[390];
   memory[97][3] = temp_mem[391];

   memory[98][0] = temp_mem[392];
   memory[98][1] = temp_mem[393];
   memory[98][2] = temp_mem[394];
   memory[98][3] = temp_mem[395];

   memory[99][0] = temp_mem[396];
   memory[99][1] = temp_mem[397];
   memory[99][2] = temp_mem[398];
   memory[99][3] = temp_mem[399];

   memory[100][0] = temp_mem[400];
   memory[100][1] = temp_mem[401];
   memory[100][2] = temp_mem[402];
   memory[100][3] = temp_mem[403];

   memory[101][0] = temp_mem[404];
   memory[101][1] = temp_mem[405];
   memory[101][2] = temp_mem[406];
   memory[101][3] = temp_mem[407];

   memory[102][0] = temp_mem[408];
   memory[102][1] = temp_mem[409];
   memory[102][2] = temp_mem[410];
   memory[102][3] = temp_mem[411];

   memory[103][0] = temp_mem[412];
   memory[103][1] = temp_mem[413];
   memory[103][2] = temp_mem[414];
   memory[103][3] = temp_mem[415];

   memory[104][0] = temp_mem[416];
   memory[104][1] = temp_mem[417];
   memory[104][2] = temp_mem[418];
   memory[104][3] = temp_mem[419];

   memory[105][0] = temp_mem[420];
   memory[105][1] = temp_mem[421];
   memory[105][2] = temp_mem[422];
   memory[105][3] = temp_mem[423];

   memory[106][0] = temp_mem[424];
   memory[106][1] = temp_mem[425];
   memory[106][2] = temp_mem[426];
   memory[106][3] = temp_mem[427];

   memory[107][0] = temp_mem[428];
   memory[107][1] = temp_mem[429];
   memory[107][2] = temp_mem[430];
   memory[107][3] = temp_mem[431];

   memory[108][0] = temp_mem[432];
   memory[108][1] = temp_mem[433];
   memory[108][2] = temp_mem[434];
   memory[108][3] = temp_mem[435];

   memory[109][0] = temp_mem[436];
   memory[109][1] = temp_mem[437];
   memory[109][2] = temp_mem[438];
   memory[109][3] = temp_mem[439];

   memory[110][0] = temp_mem[440];
   memory[110][1] = temp_mem[441];
   memory[110][2] = temp_mem[442];
   memory[110][3] = temp_mem[443];

   memory[111][0] = temp_mem[444];
   memory[111][1] = temp_mem[445];
   memory[111][2] = temp_mem[446];
   memory[111][3] = temp_mem[447];

   memory[112][0] = temp_mem[448];
   memory[112][1] = temp_mem[449];
   memory[112][2] = temp_mem[450];
   memory[112][3] = temp_mem[451];

   memory[113][0] = temp_mem[452];
   memory[113][1] = temp_mem[453];
   memory[113][2] = temp_mem[454];
   memory[113][3] = temp_mem[455];

   memory[114][0] = temp_mem[456];
   memory[114][1] = temp_mem[457];
   memory[114][2] = temp_mem[458];
   memory[114][3] = temp_mem[459];

   memory[115][0] = temp_mem[460];
   memory[115][1] = temp_mem[461];
   memory[115][2] = temp_mem[462];
   memory[115][3] = temp_mem[463];

   memory[116][0] = temp_mem[464];
   memory[116][1] = temp_mem[465];
   memory[116][2] = temp_mem[466];
   memory[116][3] = temp_mem[467];

   memory[117][0] = temp_mem[468];
   memory[117][1] = temp_mem[469];
   memory[117][2] = temp_mem[470];
   memory[117][3] = temp_mem[471];

   memory[118][0] = temp_mem[472];
   memory[118][1] = temp_mem[473];
   memory[118][2] = temp_mem[474];
   memory[118][3] = temp_mem[475];

   memory[119][0] = temp_mem[476];
   memory[119][1] = temp_mem[477];
   memory[119][2] = temp_mem[478];
   memory[119][3] = temp_mem[479];

   memory[120][0] = temp_mem[480];
   memory[120][1] = temp_mem[481];
   memory[120][2] = temp_mem[482];
   memory[120][3] = temp_mem[483];

   memory[121][0] = temp_mem[484];
   memory[121][1] = temp_mem[485];
   memory[121][2] = temp_mem[486];
   memory[121][3] = temp_mem[487];

   memory[122][0] = temp_mem[488];
   memory[122][1] = temp_mem[489];
   memory[122][2] = temp_mem[490];
   memory[122][3] = temp_mem[491];

   memory[123][0] = temp_mem[492];
   memory[123][1] = temp_mem[493];
   memory[123][2] = temp_mem[494];
   memory[123][3] = temp_mem[495];

   memory[124][0] = temp_mem[496];
   memory[124][1] = temp_mem[497];
   memory[124][2] = temp_mem[498];
   memory[124][3] = temp_mem[499];

   memory[125][0] = temp_mem[500];
   memory[125][1] = temp_mem[501];
   memory[125][2] = temp_mem[502];
   memory[125][3] = temp_mem[503];

   memory[126][0] = temp_mem[504];
   memory[126][1] = temp_mem[505];
   memory[126][2] = temp_mem[506];
   memory[126][3] = temp_mem[507];

   memory[127][0] = temp_mem[508];
   memory[127][1] = temp_mem[509];
   memory[127][2] = temp_mem[510];
   memory[127][3] = temp_mem[511];

   memory[128][0] = temp_mem[512];
   memory[128][1] = temp_mem[513];
   memory[128][2] = temp_mem[514];
   memory[128][3] = temp_mem[515];

   memory[129][0] = temp_mem[516];
   memory[129][1] = temp_mem[517];
   memory[129][2] = temp_mem[518];
   memory[129][3] = temp_mem[519];

   memory[130][0] = temp_mem[520];
   memory[130][1] = temp_mem[521];
   memory[130][2] = temp_mem[522];
   memory[130][3] = temp_mem[523];

   memory[131][0] = temp_mem[524];
   memory[131][1] = temp_mem[525];
   memory[131][2] = temp_mem[526];
   memory[131][3] = temp_mem[527];

   memory[132][0] = temp_mem[528];
   memory[132][1] = temp_mem[529];
   memory[132][2] = temp_mem[530];
   memory[132][3] = temp_mem[531];

   memory[133][0] = temp_mem[532];
   memory[133][1] = temp_mem[533];
   memory[133][2] = temp_mem[534];
   memory[133][3] = temp_mem[535];

   memory[134][0] = temp_mem[536];
   memory[134][1] = temp_mem[537];
   memory[134][2] = temp_mem[538];
   memory[134][3] = temp_mem[539];

   memory[135][0] = temp_mem[540];
   memory[135][1] = temp_mem[541];
   memory[135][2] = temp_mem[542];
   memory[135][3] = temp_mem[543];

   memory[136][0] = temp_mem[544];
   memory[136][1] = temp_mem[545];
   memory[136][2] = temp_mem[546];
   memory[136][3] = temp_mem[547];

   memory[137][0] = temp_mem[548];
   memory[137][1] = temp_mem[549];
   memory[137][2] = temp_mem[550];
   memory[137][3] = temp_mem[551];

   memory[138][0] = temp_mem[552];
   memory[138][1] = temp_mem[553];
   memory[138][2] = temp_mem[554];
   memory[138][3] = temp_mem[555];

   memory[139][0] = temp_mem[556];
   memory[139][1] = temp_mem[557];
   memory[139][2] = temp_mem[558];
   memory[139][3] = temp_mem[559];

   memory[140][0] = temp_mem[560];
   memory[140][1] = temp_mem[561];
   memory[140][2] = temp_mem[562];
   memory[140][3] = temp_mem[563];

   memory[141][0] = temp_mem[564];
   memory[141][1] = temp_mem[565];
   memory[141][2] = temp_mem[566];
   memory[141][3] = temp_mem[567];

   memory[142][0] = temp_mem[568];
   memory[142][1] = temp_mem[569];
   memory[142][2] = temp_mem[570];
   memory[142][3] = temp_mem[571];

   memory[143][0] = temp_mem[572];
   memory[143][1] = temp_mem[573];
   memory[143][2] = temp_mem[574];
   memory[143][3] = temp_mem[575];

   memory[144][0] = temp_mem[576];
   memory[144][1] = temp_mem[577];
   memory[144][2] = temp_mem[578];
   memory[144][3] = temp_mem[579];

   memory[145][0] = temp_mem[580];
   memory[145][1] = temp_mem[581];
   memory[145][2] = temp_mem[582];
   memory[145][3] = temp_mem[583];

   memory[146][0] = temp_mem[584];
   memory[146][1] = temp_mem[585];
   memory[146][2] = temp_mem[586];
   memory[146][3] = temp_mem[587];

   memory[147][0] = temp_mem[588];
   memory[147][1] = temp_mem[589];
   memory[147][2] = temp_mem[590];
   memory[147][3] = temp_mem[591];

   memory[148][0] = temp_mem[592];
   memory[148][1] = temp_mem[593];
   memory[148][2] = temp_mem[594];
   memory[148][3] = temp_mem[595];

   memory[149][0] = temp_mem[596];
   memory[149][1] = temp_mem[597];
   memory[149][2] = temp_mem[598];
   memory[149][3] = temp_mem[599];

   memory[150][0] = temp_mem[600];
   memory[150][1] = temp_mem[601];
   memory[150][2] = temp_mem[602];
   memory[150][3] = temp_mem[603];

   memory[151][0] = temp_mem[604];
   memory[151][1] = temp_mem[605];
   memory[151][2] = temp_mem[606];
   memory[151][3] = temp_mem[607];

   memory[152][0] = temp_mem[608];
   memory[152][1] = temp_mem[609];
   memory[152][2] = temp_mem[610];
   memory[152][3] = temp_mem[611];

   memory[153][0] = temp_mem[612];
   memory[153][1] = temp_mem[613];
   memory[153][2] = temp_mem[614];
   memory[153][3] = temp_mem[615];

   memory[154][0] = temp_mem[616];
   memory[154][1] = temp_mem[617];
   memory[154][2] = temp_mem[618];
   memory[154][3] = temp_mem[619];

   memory[155][0] = temp_mem[620];
   memory[155][1] = temp_mem[621];
   memory[155][2] = temp_mem[622];
   memory[155][3] = temp_mem[623];

   memory[156][0] = temp_mem[624];
   memory[156][1] = temp_mem[625];
   memory[156][2] = temp_mem[626];
   memory[156][3] = temp_mem[627];

   memory[157][0] = temp_mem[628];
   memory[157][1] = temp_mem[629];
   memory[157][2] = temp_mem[630];
   memory[157][3] = temp_mem[631];

   memory[158][0] = temp_mem[632];
   memory[158][1] = temp_mem[633];
   memory[158][2] = temp_mem[634];
   memory[158][3] = temp_mem[635];

   memory[159][0] = temp_mem[636];
   memory[159][1] = temp_mem[637];
   memory[159][2] = temp_mem[638];
   memory[159][3] = temp_mem[639];

   memory[160][0] = temp_mem[640];
   memory[160][1] = temp_mem[641];
   memory[160][2] = temp_mem[642];
   memory[160][3] = temp_mem[643];

   memory[161][0] = temp_mem[644];
   memory[161][1] = temp_mem[645];
   memory[161][2] = temp_mem[646];
   memory[161][3] = temp_mem[647];

   memory[162][0] = temp_mem[648];
   memory[162][1] = temp_mem[649];
   memory[162][2] = temp_mem[650];
   memory[162][3] = temp_mem[651];

   memory[163][0] = temp_mem[652];
   memory[163][1] = temp_mem[653];
   memory[163][2] = temp_mem[654];
   memory[163][3] = temp_mem[655];

   memory[164][0] = temp_mem[656];
   memory[164][1] = temp_mem[657];
   memory[164][2] = temp_mem[658];
   memory[164][3] = temp_mem[659];

   memory[165][0] = temp_mem[660];
   memory[165][1] = temp_mem[661];
   memory[165][2] = temp_mem[662];
   memory[165][3] = temp_mem[663];

   memory[166][0] = temp_mem[664];
   memory[166][1] = temp_mem[665];
   memory[166][2] = temp_mem[666];
   memory[166][3] = temp_mem[667];

   memory[167][0] = temp_mem[668];
   memory[167][1] = temp_mem[669];
   memory[167][2] = temp_mem[670];
   memory[167][3] = temp_mem[671];

   memory[168][0] = temp_mem[672];
   memory[168][1] = temp_mem[673];
   memory[168][2] = temp_mem[674];
   memory[168][3] = temp_mem[675];

   memory[169][0] = temp_mem[676];
   memory[169][1] = temp_mem[677];
   memory[169][2] = temp_mem[678];
   memory[169][3] = temp_mem[679];

   memory[170][0] = temp_mem[680];
   memory[170][1] = temp_mem[681];
   memory[170][2] = temp_mem[682];
   memory[170][3] = temp_mem[683];

   memory[171][0] = temp_mem[684];
   memory[171][1] = temp_mem[685];
   memory[171][2] = temp_mem[686];
   memory[171][3] = temp_mem[687];

   memory[172][0] = temp_mem[688];
   memory[172][1] = temp_mem[689];
   memory[172][2] = temp_mem[690];
   memory[172][3] = temp_mem[691];

   memory[173][0] = temp_mem[692];
   memory[173][1] = temp_mem[693];
   memory[173][2] = temp_mem[694];
   memory[173][3] = temp_mem[695];

   memory[174][0] = temp_mem[696];
   memory[174][1] = temp_mem[697];
   memory[174][2] = temp_mem[698];
   memory[174][3] = temp_mem[699];

   memory[175][0] = temp_mem[700];
   memory[175][1] = temp_mem[701];
   memory[175][2] = temp_mem[702];
   memory[175][3] = temp_mem[703];

   memory[176][0] = temp_mem[704];
   memory[176][1] = temp_mem[705];
   memory[176][2] = temp_mem[706];
   memory[176][3] = temp_mem[707];

   memory[177][0] = temp_mem[708];
   memory[177][1] = temp_mem[709];
   memory[177][2] = temp_mem[710];
   memory[177][3] = temp_mem[711];

   memory[178][0] = temp_mem[712];
   memory[178][1] = temp_mem[713];
   memory[178][2] = temp_mem[714];
   memory[178][3] = temp_mem[715];

   memory[179][0] = temp_mem[716];
   memory[179][1] = temp_mem[717];
   memory[179][2] = temp_mem[718];
   memory[179][3] = temp_mem[719];

   memory[180][0] = temp_mem[720];
   memory[180][1] = temp_mem[721];
   memory[180][2] = temp_mem[722];
   memory[180][3] = temp_mem[723];

   memory[181][0] = temp_mem[724];
   memory[181][1] = temp_mem[725];
   memory[181][2] = temp_mem[726];
   memory[181][3] = temp_mem[727];

   memory[182][0] = temp_mem[728];
   memory[182][1] = temp_mem[729];
   memory[182][2] = temp_mem[730];
   memory[182][3] = temp_mem[731];

   memory[183][0] = temp_mem[732];
   memory[183][1] = temp_mem[733];
   memory[183][2] = temp_mem[734];
   memory[183][3] = temp_mem[735];

   memory[184][0] = temp_mem[736];
   memory[184][1] = temp_mem[737];
   memory[184][2] = temp_mem[738];
   memory[184][3] = temp_mem[739];

   memory[185][0] = temp_mem[740];
   memory[185][1] = temp_mem[741];
   memory[185][2] = temp_mem[742];
   memory[185][3] = temp_mem[743];

   memory[186][0] = temp_mem[744];
   memory[186][1] = temp_mem[745];
   memory[186][2] = temp_mem[746];
   memory[186][3] = temp_mem[747];

   memory[187][0] = temp_mem[748];
   memory[187][1] = temp_mem[749];
   memory[187][2] = temp_mem[750];
   memory[187][3] = temp_mem[751];

   memory[188][0] = temp_mem[752];
   memory[188][1] = temp_mem[753];
   memory[188][2] = temp_mem[754];
   memory[188][3] = temp_mem[755];

   memory[189][0] = temp_mem[756];
   memory[189][1] = temp_mem[757];
   memory[189][2] = temp_mem[758];
   memory[189][3] = temp_mem[759];

   memory[190][0] = temp_mem[760];
   memory[190][1] = temp_mem[761];
   memory[190][2] = temp_mem[762];
   memory[190][3] = temp_mem[763];

   memory[191][0] = temp_mem[764];
   memory[191][1] = temp_mem[765];
   memory[191][2] = temp_mem[766];
   memory[191][3] = temp_mem[767];

   memory[192][0] = temp_mem[768];
   memory[192][1] = temp_mem[769];
   memory[192][2] = temp_mem[770];
   memory[192][3] = temp_mem[771];

   memory[193][0] = temp_mem[772];
   memory[193][1] = temp_mem[773];
   memory[193][2] = temp_mem[774];
   memory[193][3] = temp_mem[775];

   memory[194][0] = temp_mem[776];
   memory[194][1] = temp_mem[777];
   memory[194][2] = temp_mem[778];
   memory[194][3] = temp_mem[779];

   memory[195][0] = temp_mem[780];
   memory[195][1] = temp_mem[781];
   memory[195][2] = temp_mem[782];
   memory[195][3] = temp_mem[783];

   memory[196][0] = temp_mem[784];
   memory[196][1] = temp_mem[785];
   memory[196][2] = temp_mem[786];
   memory[196][3] = temp_mem[787];

   memory[197][0] = temp_mem[788];
   memory[197][1] = temp_mem[789];
   memory[197][2] = temp_mem[790];
   memory[197][3] = temp_mem[791];

   memory[198][0] = temp_mem[792];
   memory[198][1] = temp_mem[793];
   memory[198][2] = temp_mem[794];
   memory[198][3] = temp_mem[795];

   memory[199][0] = temp_mem[796];
   memory[199][1] = temp_mem[797];
   memory[199][2] = temp_mem[798];
   memory[199][3] = temp_mem[799];

   memory[200][0] = temp_mem[800];
   memory[200][1] = temp_mem[801];
   memory[200][2] = temp_mem[802];
   memory[200][3] = temp_mem[803];

   memory[201][0] = temp_mem[804];
   memory[201][1] = temp_mem[805];
   memory[201][2] = temp_mem[806];
   memory[201][3] = temp_mem[807];

   memory[202][0] = temp_mem[808];
   memory[202][1] = temp_mem[809];
   memory[202][2] = temp_mem[810];
   memory[202][3] = temp_mem[811];

   memory[203][0] = temp_mem[812];
   memory[203][1] = temp_mem[813];
   memory[203][2] = temp_mem[814];
   memory[203][3] = temp_mem[815];

   memory[204][0] = temp_mem[816];
   memory[204][1] = temp_mem[817];
   memory[204][2] = temp_mem[818];
   memory[204][3] = temp_mem[819];

   memory[205][0] = temp_mem[820];
   memory[205][1] = temp_mem[821];
   memory[205][2] = temp_mem[822];
   memory[205][3] = temp_mem[823];

   memory[206][0] = temp_mem[824];
   memory[206][1] = temp_mem[825];
   memory[206][2] = temp_mem[826];
   memory[206][3] = temp_mem[827];

   memory[207][0] = temp_mem[828];
   memory[207][1] = temp_mem[829];
   memory[207][2] = temp_mem[830];
   memory[207][3] = temp_mem[831];

   memory[208][0] = temp_mem[832];
   memory[208][1] = temp_mem[833];
   memory[208][2] = temp_mem[834];
   memory[208][3] = temp_mem[835];

   memory[209][0] = temp_mem[836];
   memory[209][1] = temp_mem[837];
   memory[209][2] = temp_mem[838];
   memory[209][3] = temp_mem[839];

   memory[210][0] = temp_mem[840];
   memory[210][1] = temp_mem[841];
   memory[210][2] = temp_mem[842];
   memory[210][3] = temp_mem[843];

   memory[211][0] = temp_mem[844];
   memory[211][1] = temp_mem[845];
   memory[211][2] = temp_mem[846];
   memory[211][3] = temp_mem[847];

   memory[212][0] = temp_mem[848];
   memory[212][1] = temp_mem[849];
   memory[212][2] = temp_mem[850];
   memory[212][3] = temp_mem[851];

   memory[213][0] = temp_mem[852];
   memory[213][1] = temp_mem[853];
   memory[213][2] = temp_mem[854];
   memory[213][3] = temp_mem[855];

   memory[214][0] = temp_mem[856];
   memory[214][1] = temp_mem[857];
   memory[214][2] = temp_mem[858];
   memory[214][3] = temp_mem[859];

   memory[215][0] = temp_mem[860];
   memory[215][1] = temp_mem[861];
   memory[215][2] = temp_mem[862];
   memory[215][3] = temp_mem[863];

   memory[216][0] = temp_mem[864];
   memory[216][1] = temp_mem[865];
   memory[216][2] = temp_mem[866];
   memory[216][3] = temp_mem[867];

   memory[217][0] = temp_mem[868];
   memory[217][1] = temp_mem[869];
   memory[217][2] = temp_mem[870];
   memory[217][3] = temp_mem[871];

   memory[218][0] = temp_mem[872];
   memory[218][1] = temp_mem[873];
   memory[218][2] = temp_mem[874];
   memory[218][3] = temp_mem[875];

   memory[219][0] = temp_mem[876];
   memory[219][1] = temp_mem[877];
   memory[219][2] = temp_mem[878];
   memory[219][3] = temp_mem[879];

   memory[220][0] = temp_mem[880];
   memory[220][1] = temp_mem[881];
   memory[220][2] = temp_mem[882];
   memory[220][3] = temp_mem[883];

   memory[221][0] = temp_mem[884];
   memory[221][1] = temp_mem[885];
   memory[221][2] = temp_mem[886];
   memory[221][3] = temp_mem[887];

   memory[222][0] = temp_mem[888];
   memory[222][1] = temp_mem[889];
   memory[222][2] = temp_mem[890];
   memory[222][3] = temp_mem[891];

   memory[223][0] = temp_mem[892];
   memory[223][1] = temp_mem[893];
   memory[223][2] = temp_mem[894];
   memory[223][3] = temp_mem[895];

   memory[224][0] = temp_mem[896];
   memory[224][1] = temp_mem[897];
   memory[224][2] = temp_mem[898];
   memory[224][3] = temp_mem[899];

   memory[225][0] = temp_mem[900];
   memory[225][1] = temp_mem[901];
   memory[225][2] = temp_mem[902];
   memory[225][3] = temp_mem[903];

   memory[226][0] = temp_mem[904];
   memory[226][1] = temp_mem[905];
   memory[226][2] = temp_mem[906];
   memory[226][3] = temp_mem[907];

   memory[227][0] = temp_mem[908];
   memory[227][1] = temp_mem[909];
   memory[227][2] = temp_mem[910];
   memory[227][3] = temp_mem[911];

   memory[228][0] = temp_mem[912];
   memory[228][1] = temp_mem[913];
   memory[228][2] = temp_mem[914];
   memory[228][3] = temp_mem[915];

   memory[229][0] = temp_mem[916];
   memory[229][1] = temp_mem[917];
   memory[229][2] = temp_mem[918];
   memory[229][3] = temp_mem[919];

   memory[230][0] = temp_mem[920];
   memory[230][1] = temp_mem[921];
   memory[230][2] = temp_mem[922];
   memory[230][3] = temp_mem[923];

   memory[231][0] = temp_mem[924];
   memory[231][1] = temp_mem[925];
   memory[231][2] = temp_mem[926];
   memory[231][3] = temp_mem[927];

   memory[232][0] = temp_mem[928];
   memory[232][1] = temp_mem[929];
   memory[232][2] = temp_mem[930];
   memory[232][3] = temp_mem[931];

   memory[233][0] = temp_mem[932];
   memory[233][1] = temp_mem[933];
   memory[233][2] = temp_mem[934];
   memory[233][3] = temp_mem[935];

   memory[234][0] = temp_mem[936];
   memory[234][1] = temp_mem[937];
   memory[234][2] = temp_mem[938];
   memory[234][3] = temp_mem[939];

   memory[235][0] = temp_mem[940];
   memory[235][1] = temp_mem[941];
   memory[235][2] = temp_mem[942];
   memory[235][3] = temp_mem[943];

   memory[236][0] = temp_mem[944];
   memory[236][1] = temp_mem[945];
   memory[236][2] = temp_mem[946];
   memory[236][3] = temp_mem[947];

   memory[237][0] = temp_mem[948];
   memory[237][1] = temp_mem[949];
   memory[237][2] = temp_mem[950];
   memory[237][3] = temp_mem[951];

   memory[238][0] = temp_mem[952];
   memory[238][1] = temp_mem[953];
   memory[238][2] = temp_mem[954];
   memory[238][3] = temp_mem[955];

   memory[239][0] = temp_mem[956];
   memory[239][1] = temp_mem[957];
   memory[239][2] = temp_mem[958];
   memory[239][3] = temp_mem[959];

   memory[240][0] = temp_mem[960];
   memory[240][1] = temp_mem[961];
   memory[240][2] = temp_mem[962];
   memory[240][3] = temp_mem[963];

   memory[241][0] = temp_mem[964];
   memory[241][1] = temp_mem[965];
   memory[241][2] = temp_mem[966];
   memory[241][3] = temp_mem[967];

   memory[242][0] = temp_mem[968];
   memory[242][1] = temp_mem[969];
   memory[242][2] = temp_mem[970];
   memory[242][3] = temp_mem[971];

   memory[243][0] = temp_mem[972];
   memory[243][1] = temp_mem[973];
   memory[243][2] = temp_mem[974];
   memory[243][3] = temp_mem[975];

   memory[244][0] = temp_mem[976];
   memory[244][1] = temp_mem[977];
   memory[244][2] = temp_mem[978];
   memory[244][3] = temp_mem[979];

   memory[245][0] = temp_mem[980];
   memory[245][1] = temp_mem[981];
   memory[245][2] = temp_mem[982];
   memory[245][3] = temp_mem[983];

   memory[246][0] = temp_mem[984];
   memory[246][1] = temp_mem[985];
   memory[246][2] = temp_mem[986];
   memory[246][3] = temp_mem[987];

   memory[247][0] = temp_mem[988];
   memory[247][1] = temp_mem[989];
   memory[247][2] = temp_mem[990];
   memory[247][3] = temp_mem[991];

   memory[248][0] = temp_mem[992];
   memory[248][1] = temp_mem[993];
   memory[248][2] = temp_mem[994];
   memory[248][3] = temp_mem[995];

   memory[249][0] = temp_mem[996];
   memory[249][1] = temp_mem[997];
   memory[249][2] = temp_mem[998];
   memory[249][3] = temp_mem[999];

   memory[250][0] = temp_mem[1000];
   memory[250][1] = temp_mem[1001];
   memory[250][2] = temp_mem[1002];
   memory[250][3] = temp_mem[1003];

   memory[251][0] = temp_mem[1004];
   memory[251][1] = temp_mem[1005];
   memory[251][2] = temp_mem[1006];
   memory[251][3] = temp_mem[1007];

   memory[252][0] = temp_mem[1008];
   memory[252][1] = temp_mem[1009];
   memory[252][2] = temp_mem[1010];
   memory[252][3] = temp_mem[1011];

   memory[253][0] = temp_mem[1012];
   memory[253][1] = temp_mem[1013];
   memory[253][2] = temp_mem[1014];
   memory[253][3] = temp_mem[1015];

   memory[254][0] = temp_mem[1016];
   memory[254][1] = temp_mem[1017];
   memory[254][2] = temp_mem[1018];
   memory[254][3] = temp_mem[1019];

   memory[255][0] = temp_mem[1020];
   memory[255][1] = temp_mem[1021];
   memory[255][2] = temp_mem[1022];
   memory[255][3] = temp_mem[1023];

   memory[256][0] = temp_mem[1024];
   memory[256][1] = temp_mem[1025];
   memory[256][2] = temp_mem[1026];
   memory[256][3] = temp_mem[1027];

   memory[257][0] = temp_mem[1028];
   memory[257][1] = temp_mem[1029];
   memory[257][2] = temp_mem[1030];
   memory[257][3] = temp_mem[1031];

   memory[258][0] = temp_mem[1032];
   memory[258][1] = temp_mem[1033];
   memory[258][2] = temp_mem[1034];
   memory[258][3] = temp_mem[1035];

   memory[259][0] = temp_mem[1036];
   memory[259][1] = temp_mem[1037];
   memory[259][2] = temp_mem[1038];
   memory[259][3] = temp_mem[1039];

   memory[260][0] = temp_mem[1040];
   memory[260][1] = temp_mem[1041];
   memory[260][2] = temp_mem[1042];
   memory[260][3] = temp_mem[1043];

   memory[261][0] = temp_mem[1044];
   memory[261][1] = temp_mem[1045];
   memory[261][2] = temp_mem[1046];
   memory[261][3] = temp_mem[1047];

   memory[262][0] = temp_mem[1048];
   memory[262][1] = temp_mem[1049];
   memory[262][2] = temp_mem[1050];
   memory[262][3] = temp_mem[1051];

   memory[263][0] = temp_mem[1052];
   memory[263][1] = temp_mem[1053];
   memory[263][2] = temp_mem[1054];
   memory[263][3] = temp_mem[1055];

   memory[264][0] = temp_mem[1056];
   memory[264][1] = temp_mem[1057];
   memory[264][2] = temp_mem[1058];
   memory[264][3] = temp_mem[1059];

   memory[265][0] = temp_mem[1060];
   memory[265][1] = temp_mem[1061];
   memory[265][2] = temp_mem[1062];
   memory[265][3] = temp_mem[1063];

   memory[266][0] = temp_mem[1064];
   memory[266][1] = temp_mem[1065];
   memory[266][2] = temp_mem[1066];
   memory[266][3] = temp_mem[1067];

   memory[267][0] = temp_mem[1068];
   memory[267][1] = temp_mem[1069];
   memory[267][2] = temp_mem[1070];
   memory[267][3] = temp_mem[1071];

   memory[268][0] = temp_mem[1072];
   memory[268][1] = temp_mem[1073];
   memory[268][2] = temp_mem[1074];
   memory[268][3] = temp_mem[1075];

   memory[269][0] = temp_mem[1076];
   memory[269][1] = temp_mem[1077];
   memory[269][2] = temp_mem[1078];
   memory[269][3] = temp_mem[1079];

   memory[270][0] = temp_mem[1080];
   memory[270][1] = temp_mem[1081];
   memory[270][2] = temp_mem[1082];
   memory[270][3] = temp_mem[1083];

   memory[271][0] = temp_mem[1084];
   memory[271][1] = temp_mem[1085];
   memory[271][2] = temp_mem[1086];
   memory[271][3] = temp_mem[1087];

   memory[272][0] = temp_mem[1088];
   memory[272][1] = temp_mem[1089];
   memory[272][2] = temp_mem[1090];
   memory[272][3] = temp_mem[1091];

   memory[273][0] = temp_mem[1092];
   memory[273][1] = temp_mem[1093];
   memory[273][2] = temp_mem[1094];
   memory[273][3] = temp_mem[1095];

   memory[274][0] = temp_mem[1096];
   memory[274][1] = temp_mem[1097];
   memory[274][2] = temp_mem[1098];
   memory[274][3] = temp_mem[1099];

   memory[275][0] = temp_mem[1100];
   memory[275][1] = temp_mem[1101];
   memory[275][2] = temp_mem[1102];
   memory[275][3] = temp_mem[1103];

   memory[276][0] = temp_mem[1104];
   memory[276][1] = temp_mem[1105];
   memory[276][2] = temp_mem[1106];
   memory[276][3] = temp_mem[1107];

   memory[277][0] = temp_mem[1108];
   memory[277][1] = temp_mem[1109];
   memory[277][2] = temp_mem[1110];
   memory[277][3] = temp_mem[1111];

   memory[278][0] = temp_mem[1112];
   memory[278][1] = temp_mem[1113];
   memory[278][2] = temp_mem[1114];
   memory[278][3] = temp_mem[1115];

   memory[279][0] = temp_mem[1116];
   memory[279][1] = temp_mem[1117];
   memory[279][2] = temp_mem[1118];
   memory[279][3] = temp_mem[1119];

   memory[280][0] = temp_mem[1120];
   memory[280][1] = temp_mem[1121];
   memory[280][2] = temp_mem[1122];
   memory[280][3] = temp_mem[1123];

   memory[281][0] = temp_mem[1124];
   memory[281][1] = temp_mem[1125];
   memory[281][2] = temp_mem[1126];
   memory[281][3] = temp_mem[1127];

   memory[282][0] = temp_mem[1128];
   memory[282][1] = temp_mem[1129];
   memory[282][2] = temp_mem[1130];
   memory[282][3] = temp_mem[1131];

   memory[283][0] = temp_mem[1132];
   memory[283][1] = temp_mem[1133];
   memory[283][2] = temp_mem[1134];
   memory[283][3] = temp_mem[1135];

   memory[284][0] = temp_mem[1136];
   memory[284][1] = temp_mem[1137];
   memory[284][2] = temp_mem[1138];
   memory[284][3] = temp_mem[1139];

   memory[285][0] = temp_mem[1140];
   memory[285][1] = temp_mem[1141];
   memory[285][2] = temp_mem[1142];
   memory[285][3] = temp_mem[1143];

   memory[286][0] = temp_mem[1144];
   memory[286][1] = temp_mem[1145];
   memory[286][2] = temp_mem[1146];
   memory[286][3] = temp_mem[1147];

   memory[287][0] = temp_mem[1148];
   memory[287][1] = temp_mem[1149];
   memory[287][2] = temp_mem[1150];
   memory[287][3] = temp_mem[1151];

   memory[288][0] = temp_mem[1152];
   memory[288][1] = temp_mem[1153];
   memory[288][2] = temp_mem[1154];
   memory[288][3] = temp_mem[1155];

   memory[289][0] = temp_mem[1156];
   memory[289][1] = temp_mem[1157];
   memory[289][2] = temp_mem[1158];
   memory[289][3] = temp_mem[1159];

   memory[290][0] = temp_mem[1160];
   memory[290][1] = temp_mem[1161];
   memory[290][2] = temp_mem[1162];
   memory[290][3] = temp_mem[1163];

   memory[291][0] = temp_mem[1164];
   memory[291][1] = temp_mem[1165];
   memory[291][2] = temp_mem[1166];
   memory[291][3] = temp_mem[1167];

   memory[292][0] = temp_mem[1168];
   memory[292][1] = temp_mem[1169];
   memory[292][2] = temp_mem[1170];
   memory[292][3] = temp_mem[1171];

   memory[293][0] = temp_mem[1172];
   memory[293][1] = temp_mem[1173];
   memory[293][2] = temp_mem[1174];
   memory[293][3] = temp_mem[1175];

   memory[294][0] = temp_mem[1176];
   memory[294][1] = temp_mem[1177];
   memory[294][2] = temp_mem[1178];
   memory[294][3] = temp_mem[1179];

   memory[295][0] = temp_mem[1180];
   memory[295][1] = temp_mem[1181];
   memory[295][2] = temp_mem[1182];
   memory[295][3] = temp_mem[1183];

   memory[296][0] = temp_mem[1184];
   memory[296][1] = temp_mem[1185];
   memory[296][2] = temp_mem[1186];
   memory[296][3] = temp_mem[1187];

   memory[297][0] = temp_mem[1188];
   memory[297][1] = temp_mem[1189];
   memory[297][2] = temp_mem[1190];
   memory[297][3] = temp_mem[1191];

   memory[298][0] = temp_mem[1192];
   memory[298][1] = temp_mem[1193];
   memory[298][2] = temp_mem[1194];
   memory[298][3] = temp_mem[1195];

   memory[299][0] = temp_mem[1196];
   memory[299][1] = temp_mem[1197];
   memory[299][2] = temp_mem[1198];
   memory[299][3] = temp_mem[1199];

   memory[300][0] = temp_mem[1200];
   memory[300][1] = temp_mem[1201];
   memory[300][2] = temp_mem[1202];
   memory[300][3] = temp_mem[1203];

   memory[301][0] = temp_mem[1204];
   memory[301][1] = temp_mem[1205];
   memory[301][2] = temp_mem[1206];
   memory[301][3] = temp_mem[1207];

   memory[302][0] = temp_mem[1208];
   memory[302][1] = temp_mem[1209];
   memory[302][2] = temp_mem[1210];
   memory[302][3] = temp_mem[1211];

   memory[303][0] = temp_mem[1212];
   memory[303][1] = temp_mem[1213];
   memory[303][2] = temp_mem[1214];
   memory[303][3] = temp_mem[1215];

   memory[304][0] = temp_mem[1216];
   memory[304][1] = temp_mem[1217];
   memory[304][2] = temp_mem[1218];
   memory[304][3] = temp_mem[1219];

   memory[305][0] = temp_mem[1220];
   memory[305][1] = temp_mem[1221];
   memory[305][2] = temp_mem[1222];
   memory[305][3] = temp_mem[1223];

   memory[306][0] = temp_mem[1224];
   memory[306][1] = temp_mem[1225];
   memory[306][2] = temp_mem[1226];
   memory[306][3] = temp_mem[1227];

   memory[307][0] = temp_mem[1228];
   memory[307][1] = temp_mem[1229];
   memory[307][2] = temp_mem[1230];
   memory[307][3] = temp_mem[1231];

   memory[308][0] = temp_mem[1232];
   memory[308][1] = temp_mem[1233];
   memory[308][2] = temp_mem[1234];
   memory[308][3] = temp_mem[1235];

   memory[309][0] = temp_mem[1236];
   memory[309][1] = temp_mem[1237];
   memory[309][2] = temp_mem[1238];
   memory[309][3] = temp_mem[1239];

   memory[310][0] = temp_mem[1240];
   memory[310][1] = temp_mem[1241];
   memory[310][2] = temp_mem[1242];
   memory[310][3] = temp_mem[1243];

   memory[311][0] = temp_mem[1244];
   memory[311][1] = temp_mem[1245];
   memory[311][2] = temp_mem[1246];
   memory[311][3] = temp_mem[1247];

   memory[312][0] = temp_mem[1248];
   memory[312][1] = temp_mem[1249];
   memory[312][2] = temp_mem[1250];
   memory[312][3] = temp_mem[1251];

   memory[313][0] = temp_mem[1252];
   memory[313][1] = temp_mem[1253];
   memory[313][2] = temp_mem[1254];
   memory[313][3] = temp_mem[1255];

   memory[314][0] = temp_mem[1256];
   memory[314][1] = temp_mem[1257];
   memory[314][2] = temp_mem[1258];
   memory[314][3] = temp_mem[1259];

   memory[315][0] = temp_mem[1260];
   memory[315][1] = temp_mem[1261];
   memory[315][2] = temp_mem[1262];
   memory[315][3] = temp_mem[1263];

   memory[316][0] = temp_mem[1264];
   memory[316][1] = temp_mem[1265];
   memory[316][2] = temp_mem[1266];
   memory[316][3] = temp_mem[1267];

   memory[317][0] = temp_mem[1268];
   memory[317][1] = temp_mem[1269];
   memory[317][2] = temp_mem[1270];
   memory[317][3] = temp_mem[1271];

   memory[318][0] = temp_mem[1272];
   memory[318][1] = temp_mem[1273];
   memory[318][2] = temp_mem[1274];
   memory[318][3] = temp_mem[1275];

   memory[319][0] = temp_mem[1276];
   memory[319][1] = temp_mem[1277];
   memory[319][2] = temp_mem[1278];
   memory[319][3] = temp_mem[1279];

   memory[320][0] = temp_mem[1280];
   memory[320][1] = temp_mem[1281];
   memory[320][2] = temp_mem[1282];
   memory[320][3] = temp_mem[1283];

   memory[321][0] = temp_mem[1284];
   memory[321][1] = temp_mem[1285];
   memory[321][2] = temp_mem[1286];
   memory[321][3] = temp_mem[1287];

   memory[322][0] = temp_mem[1288];
   memory[322][1] = temp_mem[1289];
   memory[322][2] = temp_mem[1290];
   memory[322][3] = temp_mem[1291];

   memory[323][0] = temp_mem[1292];
   memory[323][1] = temp_mem[1293];
   memory[323][2] = temp_mem[1294];
   memory[323][3] = temp_mem[1295];

   memory[324][0] = temp_mem[1296];
   memory[324][1] = temp_mem[1297];
   memory[324][2] = temp_mem[1298];
   memory[324][3] = temp_mem[1299];

   memory[325][0] = temp_mem[1300];
   memory[325][1] = temp_mem[1301];
   memory[325][2] = temp_mem[1302];
   memory[325][3] = temp_mem[1303];

   memory[326][0] = temp_mem[1304];
   memory[326][1] = temp_mem[1305];
   memory[326][2] = temp_mem[1306];
   memory[326][3] = temp_mem[1307];

   memory[327][0] = temp_mem[1308];
   memory[327][1] = temp_mem[1309];
   memory[327][2] = temp_mem[1310];
   memory[327][3] = temp_mem[1311];

   memory[328][0] = temp_mem[1312];
   memory[328][1] = temp_mem[1313];
   memory[328][2] = temp_mem[1314];
   memory[328][3] = temp_mem[1315];

   memory[329][0] = temp_mem[1316];
   memory[329][1] = temp_mem[1317];
   memory[329][2] = temp_mem[1318];
   memory[329][3] = temp_mem[1319];

   memory[330][0] = temp_mem[1320];
   memory[330][1] = temp_mem[1321];
   memory[330][2] = temp_mem[1322];
   memory[330][3] = temp_mem[1323];

   memory[331][0] = temp_mem[1324];
   memory[331][1] = temp_mem[1325];
   memory[331][2] = temp_mem[1326];
   memory[331][3] = temp_mem[1327];

   memory[332][0] = temp_mem[1328];
   memory[332][1] = temp_mem[1329];
   memory[332][2] = temp_mem[1330];
   memory[332][3] = temp_mem[1331];

   memory[333][0] = temp_mem[1332];
   memory[333][1] = temp_mem[1333];
   memory[333][2] = temp_mem[1334];
   memory[333][3] = temp_mem[1335];

   memory[334][0] = temp_mem[1336];
   memory[334][1] = temp_mem[1337];
   memory[334][2] = temp_mem[1338];
   memory[334][3] = temp_mem[1339];

   memory[335][0] = temp_mem[1340];
   memory[335][1] = temp_mem[1341];
   memory[335][2] = temp_mem[1342];
   memory[335][3] = temp_mem[1343];

   memory[336][0] = temp_mem[1344];
   memory[336][1] = temp_mem[1345];
   memory[336][2] = temp_mem[1346];
   memory[336][3] = temp_mem[1347];

   memory[337][0] = temp_mem[1348];
   memory[337][1] = temp_mem[1349];
   memory[337][2] = temp_mem[1350];
   memory[337][3] = temp_mem[1351];

   memory[338][0] = temp_mem[1352];
   memory[338][1] = temp_mem[1353];
   memory[338][2] = temp_mem[1354];
   memory[338][3] = temp_mem[1355];

   memory[339][0] = temp_mem[1356];
   memory[339][1] = temp_mem[1357];
   memory[339][2] = temp_mem[1358];
   memory[339][3] = temp_mem[1359];

   memory[340][0] = temp_mem[1360];
   memory[340][1] = temp_mem[1361];
   memory[340][2] = temp_mem[1362];
   memory[340][3] = temp_mem[1363];

   memory[341][0] = temp_mem[1364];
   memory[341][1] = temp_mem[1365];
   memory[341][2] = temp_mem[1366];
   memory[341][3] = temp_mem[1367];

   memory[342][0] = temp_mem[1368];
   memory[342][1] = temp_mem[1369];
   memory[342][2] = temp_mem[1370];
   memory[342][3] = temp_mem[1371];

   memory[343][0] = temp_mem[1372];
   memory[343][1] = temp_mem[1373];
   memory[343][2] = temp_mem[1374];
   memory[343][3] = temp_mem[1375];

   memory[344][0] = temp_mem[1376];
   memory[344][1] = temp_mem[1377];
   memory[344][2] = temp_mem[1378];
   memory[344][3] = temp_mem[1379];

   memory[345][0] = temp_mem[1380];
   memory[345][1] = temp_mem[1381];
   memory[345][2] = temp_mem[1382];
   memory[345][3] = temp_mem[1383];

   memory[346][0] = temp_mem[1384];
   memory[346][1] = temp_mem[1385];
   memory[346][2] = temp_mem[1386];
   memory[346][3] = temp_mem[1387];

   memory[347][0] = temp_mem[1388];
   memory[347][1] = temp_mem[1389];
   memory[347][2] = temp_mem[1390];
   memory[347][3] = temp_mem[1391];

   memory[348][0] = temp_mem[1392];
   memory[348][1] = temp_mem[1393];
   memory[348][2] = temp_mem[1394];
   memory[348][3] = temp_mem[1395];

   memory[349][0] = temp_mem[1396];
   memory[349][1] = temp_mem[1397];
   memory[349][2] = temp_mem[1398];
   memory[349][3] = temp_mem[1399];

   memory[350][0] = temp_mem[1400];
   memory[350][1] = temp_mem[1401];
   memory[350][2] = temp_mem[1402];
   memory[350][3] = temp_mem[1403];

   memory[351][0] = temp_mem[1404];
   memory[351][1] = temp_mem[1405];
   memory[351][2] = temp_mem[1406];
   memory[351][3] = temp_mem[1407];

   memory[352][0] = temp_mem[1408];
   memory[352][1] = temp_mem[1409];
   memory[352][2] = temp_mem[1410];
   memory[352][3] = temp_mem[1411];

   memory[353][0] = temp_mem[1412];
   memory[353][1] = temp_mem[1413];
   memory[353][2] = temp_mem[1414];
   memory[353][3] = temp_mem[1415];

   memory[354][0] = temp_mem[1416];
   memory[354][1] = temp_mem[1417];
   memory[354][2] = temp_mem[1418];
   memory[354][3] = temp_mem[1419];

   memory[355][0] = temp_mem[1420];
   memory[355][1] = temp_mem[1421];
   memory[355][2] = temp_mem[1422];
   memory[355][3] = temp_mem[1423];

   memory[356][0] = temp_mem[1424];
   memory[356][1] = temp_mem[1425];
   memory[356][2] = temp_mem[1426];
   memory[356][3] = temp_mem[1427];

   memory[357][0] = temp_mem[1428];
   memory[357][1] = temp_mem[1429];
   memory[357][2] = temp_mem[1430];
   memory[357][3] = temp_mem[1431];

   memory[358][0] = temp_mem[1432];
   memory[358][1] = temp_mem[1433];
   memory[358][2] = temp_mem[1434];
   memory[358][3] = temp_mem[1435];

   memory[359][0] = temp_mem[1436];
   memory[359][1] = temp_mem[1437];
   memory[359][2] = temp_mem[1438];
   memory[359][3] = temp_mem[1439];

   memory[360][0] = temp_mem[1440];
   memory[360][1] = temp_mem[1441];
   memory[360][2] = temp_mem[1442];
   memory[360][3] = temp_mem[1443];

   memory[361][0] = temp_mem[1444];
   memory[361][1] = temp_mem[1445];
   memory[361][2] = temp_mem[1446];
   memory[361][3] = temp_mem[1447];

   memory[362][0] = temp_mem[1448];
   memory[362][1] = temp_mem[1449];
   memory[362][2] = temp_mem[1450];
   memory[362][3] = temp_mem[1451];

   memory[363][0] = temp_mem[1452];
   memory[363][1] = temp_mem[1453];
   memory[363][2] = temp_mem[1454];
   memory[363][3] = temp_mem[1455];

   memory[364][0] = temp_mem[1456];
   memory[364][1] = temp_mem[1457];
   memory[364][2] = temp_mem[1458];
   memory[364][3] = temp_mem[1459];

   memory[365][0] = temp_mem[1460];
   memory[365][1] = temp_mem[1461];
   memory[365][2] = temp_mem[1462];
   memory[365][3] = temp_mem[1463];

   memory[366][0] = temp_mem[1464];
   memory[366][1] = temp_mem[1465];
   memory[366][2] = temp_mem[1466];
   memory[366][3] = temp_mem[1467];

   memory[367][0] = temp_mem[1468];
   memory[367][1] = temp_mem[1469];
   memory[367][2] = temp_mem[1470];
   memory[367][3] = temp_mem[1471];

   memory[368][0] = temp_mem[1472];
   memory[368][1] = temp_mem[1473];
   memory[368][2] = temp_mem[1474];
   memory[368][3] = temp_mem[1475];

   memory[369][0] = temp_mem[1476];
   memory[369][1] = temp_mem[1477];
   memory[369][2] = temp_mem[1478];
   memory[369][3] = temp_mem[1479];

   memory[370][0] = temp_mem[1480];
   memory[370][1] = temp_mem[1481];
   memory[370][2] = temp_mem[1482];
   memory[370][3] = temp_mem[1483];

   memory[371][0] = temp_mem[1484];
   memory[371][1] = temp_mem[1485];
   memory[371][2] = temp_mem[1486];
   memory[371][3] = temp_mem[1487];

   memory[372][0] = temp_mem[1488];
   memory[372][1] = temp_mem[1489];
   memory[372][2] = temp_mem[1490];
   memory[372][3] = temp_mem[1491];

   memory[373][0] = temp_mem[1492];
   memory[373][1] = temp_mem[1493];
   memory[373][2] = temp_mem[1494];
   memory[373][3] = temp_mem[1495];

   memory[374][0] = temp_mem[1496];
   memory[374][1] = temp_mem[1497];
   memory[374][2] = temp_mem[1498];
   memory[374][3] = temp_mem[1499];

   memory[375][0] = temp_mem[1500];
   memory[375][1] = temp_mem[1501];
   memory[375][2] = temp_mem[1502];
   memory[375][3] = temp_mem[1503];

   memory[376][0] = temp_mem[1504];
   memory[376][1] = temp_mem[1505];
   memory[376][2] = temp_mem[1506];
   memory[376][3] = temp_mem[1507];

   memory[377][0] = temp_mem[1508];
   memory[377][1] = temp_mem[1509];
   memory[377][2] = temp_mem[1510];
   memory[377][3] = temp_mem[1511];

   memory[378][0] = temp_mem[1512];
   memory[378][1] = temp_mem[1513];
   memory[378][2] = temp_mem[1514];
   memory[378][3] = temp_mem[1515];

   memory[379][0] = temp_mem[1516];
   memory[379][1] = temp_mem[1517];
   memory[379][2] = temp_mem[1518];
   memory[379][3] = temp_mem[1519];

   memory[380][0] = temp_mem[1520];
   memory[380][1] = temp_mem[1521];
   memory[380][2] = temp_mem[1522];
   memory[380][3] = temp_mem[1523];

   memory[381][0] = temp_mem[1524];
   memory[381][1] = temp_mem[1525];
   memory[381][2] = temp_mem[1526];
   memory[381][3] = temp_mem[1527];

   memory[382][0] = temp_mem[1528];
   memory[382][1] = temp_mem[1529];
   memory[382][2] = temp_mem[1530];
   memory[382][3] = temp_mem[1531];

   memory[383][0] = temp_mem[1532];
   memory[383][1] = temp_mem[1533];
   memory[383][2] = temp_mem[1534];
   memory[383][3] = temp_mem[1535];

   memory[384][0] = temp_mem[1536];
   memory[384][1] = temp_mem[1537];
   memory[384][2] = temp_mem[1538];
   memory[384][3] = temp_mem[1539];

   memory[385][0] = temp_mem[1540];
   memory[385][1] = temp_mem[1541];
   memory[385][2] = temp_mem[1542];
   memory[385][3] = temp_mem[1543];

   memory[386][0] = temp_mem[1544];
   memory[386][1] = temp_mem[1545];
   memory[386][2] = temp_mem[1546];
   memory[386][3] = temp_mem[1547];

   memory[387][0] = temp_mem[1548];
   memory[387][1] = temp_mem[1549];
   memory[387][2] = temp_mem[1550];
   memory[387][3] = temp_mem[1551];

   memory[388][0] = temp_mem[1552];
   memory[388][1] = temp_mem[1553];
   memory[388][2] = temp_mem[1554];
   memory[388][3] = temp_mem[1555];

   memory[389][0] = temp_mem[1556];
   memory[389][1] = temp_mem[1557];
   memory[389][2] = temp_mem[1558];
   memory[389][3] = temp_mem[1559];

   memory[390][0] = temp_mem[1560];
   memory[390][1] = temp_mem[1561];
   memory[390][2] = temp_mem[1562];
   memory[390][3] = temp_mem[1563];

   memory[391][0] = temp_mem[1564];
   memory[391][1] = temp_mem[1565];
   memory[391][2] = temp_mem[1566];
   memory[391][3] = temp_mem[1567];

   memory[392][0] = temp_mem[1568];
   memory[392][1] = temp_mem[1569];
   memory[392][2] = temp_mem[1570];
   memory[392][3] = temp_mem[1571];

   memory[393][0] = temp_mem[1572];
   memory[393][1] = temp_mem[1573];
   memory[393][2] = temp_mem[1574];
   memory[393][3] = temp_mem[1575];

   memory[394][0] = temp_mem[1576];
   memory[394][1] = temp_mem[1577];
   memory[394][2] = temp_mem[1578];
   memory[394][3] = temp_mem[1579];

   memory[395][0] = temp_mem[1580];
   memory[395][1] = temp_mem[1581];
   memory[395][2] = temp_mem[1582];
   memory[395][3] = temp_mem[1583];

   memory[396][0] = temp_mem[1584];
   memory[396][1] = temp_mem[1585];
   memory[396][2] = temp_mem[1586];
   memory[396][3] = temp_mem[1587];

   memory[397][0] = temp_mem[1588];
   memory[397][1] = temp_mem[1589];
   memory[397][2] = temp_mem[1590];
   memory[397][3] = temp_mem[1591];

   memory[398][0] = temp_mem[1592];
   memory[398][1] = temp_mem[1593];
   memory[398][2] = temp_mem[1594];
   memory[398][3] = temp_mem[1595];

   memory[399][0] = temp_mem[1596];
   memory[399][1] = temp_mem[1597];
   memory[399][2] = temp_mem[1598];
   memory[399][3] = temp_mem[1599];

   memory[400][0] = temp_mem[1600];
   memory[400][1] = temp_mem[1601];
   memory[400][2] = temp_mem[1602];
   memory[400][3] = temp_mem[1603];

   memory[401][0] = temp_mem[1604];
   memory[401][1] = temp_mem[1605];
   memory[401][2] = temp_mem[1606];
   memory[401][3] = temp_mem[1607];

   memory[402][0] = temp_mem[1608];
   memory[402][1] = temp_mem[1609];
   memory[402][2] = temp_mem[1610];
   memory[402][3] = temp_mem[1611];

   memory[403][0] = temp_mem[1612];
   memory[403][1] = temp_mem[1613];
   memory[403][2] = temp_mem[1614];
   memory[403][3] = temp_mem[1615];

   memory[404][0] = temp_mem[1616];
   memory[404][1] = temp_mem[1617];
   memory[404][2] = temp_mem[1618];
   memory[404][3] = temp_mem[1619];

   memory[405][0] = temp_mem[1620];
   memory[405][1] = temp_mem[1621];
   memory[405][2] = temp_mem[1622];
   memory[405][3] = temp_mem[1623];

   memory[406][0] = temp_mem[1624];
   memory[406][1] = temp_mem[1625];
   memory[406][2] = temp_mem[1626];
   memory[406][3] = temp_mem[1627];

   memory[407][0] = temp_mem[1628];
   memory[407][1] = temp_mem[1629];
   memory[407][2] = temp_mem[1630];
   memory[407][3] = temp_mem[1631];

   memory[408][0] = temp_mem[1632];
   memory[408][1] = temp_mem[1633];
   memory[408][2] = temp_mem[1634];
   memory[408][3] = temp_mem[1635];

   memory[409][0] = temp_mem[1636];
   memory[409][1] = temp_mem[1637];
   memory[409][2] = temp_mem[1638];
   memory[409][3] = temp_mem[1639];

   memory[410][0] = temp_mem[1640];
   memory[410][1] = temp_mem[1641];
   memory[410][2] = temp_mem[1642];
   memory[410][3] = temp_mem[1643];

   memory[411][0] = temp_mem[1644];
   memory[411][1] = temp_mem[1645];
   memory[411][2] = temp_mem[1646];
   memory[411][3] = temp_mem[1647];

   memory[412][0] = temp_mem[1648];
   memory[412][1] = temp_mem[1649];
   memory[412][2] = temp_mem[1650];
   memory[412][3] = temp_mem[1651];

   memory[413][0] = temp_mem[1652];
   memory[413][1] = temp_mem[1653];
   memory[413][2] = temp_mem[1654];
   memory[413][3] = temp_mem[1655];

   memory[414][0] = temp_mem[1656];
   memory[414][1] = temp_mem[1657];
   memory[414][2] = temp_mem[1658];
   memory[414][3] = temp_mem[1659];

   memory[415][0] = temp_mem[1660];
   memory[415][1] = temp_mem[1661];
   memory[415][2] = temp_mem[1662];
   memory[415][3] = temp_mem[1663];

   memory[416][0] = temp_mem[1664];
   memory[416][1] = temp_mem[1665];
   memory[416][2] = temp_mem[1666];
   memory[416][3] = temp_mem[1667];

   memory[417][0] = temp_mem[1668];
   memory[417][1] = temp_mem[1669];
   memory[417][2] = temp_mem[1670];
   memory[417][3] = temp_mem[1671];

   memory[418][0] = temp_mem[1672];
   memory[418][1] = temp_mem[1673];
   memory[418][2] = temp_mem[1674];
   memory[418][3] = temp_mem[1675];

   memory[419][0] = temp_mem[1676];
   memory[419][1] = temp_mem[1677];
   memory[419][2] = temp_mem[1678];
   memory[419][3] = temp_mem[1679];

   memory[420][0] = temp_mem[1680];
   memory[420][1] = temp_mem[1681];
   memory[420][2] = temp_mem[1682];
   memory[420][3] = temp_mem[1683];

   memory[421][0] = temp_mem[1684];
   memory[421][1] = temp_mem[1685];
   memory[421][2] = temp_mem[1686];
   memory[421][3] = temp_mem[1687];

   memory[422][0] = temp_mem[1688];
   memory[422][1] = temp_mem[1689];
   memory[422][2] = temp_mem[1690];
   memory[422][3] = temp_mem[1691];

   memory[423][0] = temp_mem[1692];
   memory[423][1] = temp_mem[1693];
   memory[423][2] = temp_mem[1694];
   memory[423][3] = temp_mem[1695];

   memory[424][0] = temp_mem[1696];
   memory[424][1] = temp_mem[1697];
   memory[424][2] = temp_mem[1698];
   memory[424][3] = temp_mem[1699];

   memory[425][0] = temp_mem[1700];
   memory[425][1] = temp_mem[1701];
   memory[425][2] = temp_mem[1702];
   memory[425][3] = temp_mem[1703];

   memory[426][0] = temp_mem[1704];
   memory[426][1] = temp_mem[1705];
   memory[426][2] = temp_mem[1706];
   memory[426][3] = temp_mem[1707];

   memory[427][0] = temp_mem[1708];
   memory[427][1] = temp_mem[1709];
   memory[427][2] = temp_mem[1710];
   memory[427][3] = temp_mem[1711];

   memory[428][0] = temp_mem[1712];
   memory[428][1] = temp_mem[1713];
   memory[428][2] = temp_mem[1714];
   memory[428][3] = temp_mem[1715];

   memory[429][0] = temp_mem[1716];
   memory[429][1] = temp_mem[1717];
   memory[429][2] = temp_mem[1718];
   memory[429][3] = temp_mem[1719];

   memory[430][0] = temp_mem[1720];
   memory[430][1] = temp_mem[1721];
   memory[430][2] = temp_mem[1722];
   memory[430][3] = temp_mem[1723];

   memory[431][0] = temp_mem[1724];
   memory[431][1] = temp_mem[1725];
   memory[431][2] = temp_mem[1726];
   memory[431][3] = temp_mem[1727];

   memory[432][0] = temp_mem[1728];
   memory[432][1] = temp_mem[1729];
   memory[432][2] = temp_mem[1730];
   memory[432][3] = temp_mem[1731];

   memory[433][0] = temp_mem[1732];
   memory[433][1] = temp_mem[1733];
   memory[433][2] = temp_mem[1734];
   memory[433][3] = temp_mem[1735];

   memory[434][0] = temp_mem[1736];
   memory[434][1] = temp_mem[1737];
   memory[434][2] = temp_mem[1738];
   memory[434][3] = temp_mem[1739];

   memory[435][0] = temp_mem[1740];
   memory[435][1] = temp_mem[1741];
   memory[435][2] = temp_mem[1742];
   memory[435][3] = temp_mem[1743];

   memory[436][0] = temp_mem[1744];
   memory[436][1] = temp_mem[1745];
   memory[436][2] = temp_mem[1746];
   memory[436][3] = temp_mem[1747];

   memory[437][0] = temp_mem[1748];
   memory[437][1] = temp_mem[1749];
   memory[437][2] = temp_mem[1750];
   memory[437][3] = temp_mem[1751];

   memory[438][0] = temp_mem[1752];
   memory[438][1] = temp_mem[1753];
   memory[438][2] = temp_mem[1754];
   memory[438][3] = temp_mem[1755];

   memory[439][0] = temp_mem[1756];
   memory[439][1] = temp_mem[1757];
   memory[439][2] = temp_mem[1758];
   memory[439][3] = temp_mem[1759];

   memory[440][0] = temp_mem[1760];
   memory[440][1] = temp_mem[1761];
   memory[440][2] = temp_mem[1762];
   memory[440][3] = temp_mem[1763];

   memory[441][0] = temp_mem[1764];
   memory[441][1] = temp_mem[1765];
   memory[441][2] = temp_mem[1766];
   memory[441][3] = temp_mem[1767];

   memory[442][0] = temp_mem[1768];
   memory[442][1] = temp_mem[1769];
   memory[442][2] = temp_mem[1770];
   memory[442][3] = temp_mem[1771];

   memory[443][0] = temp_mem[1772];
   memory[443][1] = temp_mem[1773];
   memory[443][2] = temp_mem[1774];
   memory[443][3] = temp_mem[1775];

   memory[444][0] = temp_mem[1776];
   memory[444][1] = temp_mem[1777];
   memory[444][2] = temp_mem[1778];
   memory[444][3] = temp_mem[1779];

   memory[445][0] = temp_mem[1780];
   memory[445][1] = temp_mem[1781];
   memory[445][2] = temp_mem[1782];
   memory[445][3] = temp_mem[1783];

   memory[446][0] = temp_mem[1784];
   memory[446][1] = temp_mem[1785];
   memory[446][2] = temp_mem[1786];
   memory[446][3] = temp_mem[1787];

   memory[447][0] = temp_mem[1788];
   memory[447][1] = temp_mem[1789];
   memory[447][2] = temp_mem[1790];
   memory[447][3] = temp_mem[1791];

   memory[448][0] = temp_mem[1792];
   memory[448][1] = temp_mem[1793];
   memory[448][2] = temp_mem[1794];
   memory[448][3] = temp_mem[1795];

   memory[449][0] = temp_mem[1796];
   memory[449][1] = temp_mem[1797];
   memory[449][2] = temp_mem[1798];
   memory[449][3] = temp_mem[1799];

   memory[450][0] = temp_mem[1800];
   memory[450][1] = temp_mem[1801];
   memory[450][2] = temp_mem[1802];
   memory[450][3] = temp_mem[1803];

   memory[451][0] = temp_mem[1804];
   memory[451][1] = temp_mem[1805];
   memory[451][2] = temp_mem[1806];
   memory[451][3] = temp_mem[1807];

   memory[452][0] = temp_mem[1808];
   memory[452][1] = temp_mem[1809];
   memory[452][2] = temp_mem[1810];
   memory[452][3] = temp_mem[1811];

   memory[453][0] = temp_mem[1812];
   memory[453][1] = temp_mem[1813];
   memory[453][2] = temp_mem[1814];
   memory[453][3] = temp_mem[1815];

   memory[454][0] = temp_mem[1816];
   memory[454][1] = temp_mem[1817];
   memory[454][2] = temp_mem[1818];
   memory[454][3] = temp_mem[1819];

   memory[455][0] = temp_mem[1820];
   memory[455][1] = temp_mem[1821];
   memory[455][2] = temp_mem[1822];
   memory[455][3] = temp_mem[1823];

   memory[456][0] = temp_mem[1824];
   memory[456][1] = temp_mem[1825];
   memory[456][2] = temp_mem[1826];
   memory[456][3] = temp_mem[1827];

   memory[457][0] = temp_mem[1828];
   memory[457][1] = temp_mem[1829];
   memory[457][2] = temp_mem[1830];
   memory[457][3] = temp_mem[1831];

   memory[458][0] = temp_mem[1832];
   memory[458][1] = temp_mem[1833];
   memory[458][2] = temp_mem[1834];
   memory[458][3] = temp_mem[1835];

   memory[459][0] = temp_mem[1836];
   memory[459][1] = temp_mem[1837];
   memory[459][2] = temp_mem[1838];
   memory[459][3] = temp_mem[1839];

   memory[460][0] = temp_mem[1840];
   memory[460][1] = temp_mem[1841];
   memory[460][2] = temp_mem[1842];
   memory[460][3] = temp_mem[1843];

   memory[461][0] = temp_mem[1844];
   memory[461][1] = temp_mem[1845];
   memory[461][2] = temp_mem[1846];
   memory[461][3] = temp_mem[1847];

   memory[462][0] = temp_mem[1848];
   memory[462][1] = temp_mem[1849];
   memory[462][2] = temp_mem[1850];
   memory[462][3] = temp_mem[1851];

   memory[463][0] = temp_mem[1852];
   memory[463][1] = temp_mem[1853];
   memory[463][2] = temp_mem[1854];
   memory[463][3] = temp_mem[1855];

   memory[464][0] = temp_mem[1856];
   memory[464][1] = temp_mem[1857];
   memory[464][2] = temp_mem[1858];
   memory[464][3] = temp_mem[1859];

   memory[465][0] = temp_mem[1860];
   memory[465][1] = temp_mem[1861];
   memory[465][2] = temp_mem[1862];
   memory[465][3] = temp_mem[1863];

   memory[466][0] = temp_mem[1864];
   memory[466][1] = temp_mem[1865];
   memory[466][2] = temp_mem[1866];
   memory[466][3] = temp_mem[1867];

   memory[467][0] = temp_mem[1868];
   memory[467][1] = temp_mem[1869];
   memory[467][2] = temp_mem[1870];
   memory[467][3] = temp_mem[1871];

   memory[468][0] = temp_mem[1872];
   memory[468][1] = temp_mem[1873];
   memory[468][2] = temp_mem[1874];
   memory[468][3] = temp_mem[1875];

   memory[469][0] = temp_mem[1876];
   memory[469][1] = temp_mem[1877];
   memory[469][2] = temp_mem[1878];
   memory[469][3] = temp_mem[1879];

   memory[470][0] = temp_mem[1880];
   memory[470][1] = temp_mem[1881];
   memory[470][2] = temp_mem[1882];
   memory[470][3] = temp_mem[1883];

   memory[471][0] = temp_mem[1884];
   memory[471][1] = temp_mem[1885];
   memory[471][2] = temp_mem[1886];
   memory[471][3] = temp_mem[1887];

   memory[472][0] = temp_mem[1888];
   memory[472][1] = temp_mem[1889];
   memory[472][2] = temp_mem[1890];
   memory[472][3] = temp_mem[1891];

   memory[473][0] = temp_mem[1892];
   memory[473][1] = temp_mem[1893];
   memory[473][2] = temp_mem[1894];
   memory[473][3] = temp_mem[1895];

   memory[474][0] = temp_mem[1896];
   memory[474][1] = temp_mem[1897];
   memory[474][2] = temp_mem[1898];
   memory[474][3] = temp_mem[1899];

   memory[475][0] = temp_mem[1900];
   memory[475][1] = temp_mem[1901];
   memory[475][2] = temp_mem[1902];
   memory[475][3] = temp_mem[1903];

   memory[476][0] = temp_mem[1904];
   memory[476][1] = temp_mem[1905];
   memory[476][2] = temp_mem[1906];
   memory[476][3] = temp_mem[1907];

   memory[477][0] = temp_mem[1908];
   memory[477][1] = temp_mem[1909];
   memory[477][2] = temp_mem[1910];
   memory[477][3] = temp_mem[1911];

   memory[478][0] = temp_mem[1912];
   memory[478][1] = temp_mem[1913];
   memory[478][2] = temp_mem[1914];
   memory[478][3] = temp_mem[1915];

   memory[479][0] = temp_mem[1916];
   memory[479][1] = temp_mem[1917];
   memory[479][2] = temp_mem[1918];
   memory[479][3] = temp_mem[1919];

   memory[480][0] = temp_mem[1920];
   memory[480][1] = temp_mem[1921];
   memory[480][2] = temp_mem[1922];
   memory[480][3] = temp_mem[1923];

   memory[481][0] = temp_mem[1924];
   memory[481][1] = temp_mem[1925];
   memory[481][2] = temp_mem[1926];
   memory[481][3] = temp_mem[1927];

   memory[482][0] = temp_mem[1928];
   memory[482][1] = temp_mem[1929];
   memory[482][2] = temp_mem[1930];
   memory[482][3] = temp_mem[1931];

   memory[483][0] = temp_mem[1932];
   memory[483][1] = temp_mem[1933];
   memory[483][2] = temp_mem[1934];
   memory[483][3] = temp_mem[1935];

   memory[484][0] = temp_mem[1936];
   memory[484][1] = temp_mem[1937];
   memory[484][2] = temp_mem[1938];
   memory[484][3] = temp_mem[1939];

   memory[485][0] = temp_mem[1940];
   memory[485][1] = temp_mem[1941];
   memory[485][2] = temp_mem[1942];
   memory[485][3] = temp_mem[1943];

   memory[486][0] = temp_mem[1944];
   memory[486][1] = temp_mem[1945];
   memory[486][2] = temp_mem[1946];
   memory[486][3] = temp_mem[1947];

   memory[487][0] = temp_mem[1948];
   memory[487][1] = temp_mem[1949];
   memory[487][2] = temp_mem[1950];
   memory[487][3] = temp_mem[1951];

   memory[488][0] = temp_mem[1952];
   memory[488][1] = temp_mem[1953];
   memory[488][2] = temp_mem[1954];
   memory[488][3] = temp_mem[1955];

   memory[489][0] = temp_mem[1956];
   memory[489][1] = temp_mem[1957];
   memory[489][2] = temp_mem[1958];
   memory[489][3] = temp_mem[1959];

   memory[490][0] = temp_mem[1960];
   memory[490][1] = temp_mem[1961];
   memory[490][2] = temp_mem[1962];
   memory[490][3] = temp_mem[1963];

   memory[491][0] = temp_mem[1964];
   memory[491][1] = temp_mem[1965];
   memory[491][2] = temp_mem[1966];
   memory[491][3] = temp_mem[1967];

   memory[492][0] = temp_mem[1968];
   memory[492][1] = temp_mem[1969];
   memory[492][2] = temp_mem[1970];
   memory[492][3] = temp_mem[1971];

   memory[493][0] = temp_mem[1972];
   memory[493][1] = temp_mem[1973];
   memory[493][2] = temp_mem[1974];
   memory[493][3] = temp_mem[1975];

   memory[494][0] = temp_mem[1976];
   memory[494][1] = temp_mem[1977];
   memory[494][2] = temp_mem[1978];
   memory[494][3] = temp_mem[1979];

   memory[495][0] = temp_mem[1980];
   memory[495][1] = temp_mem[1981];
   memory[495][2] = temp_mem[1982];
   memory[495][3] = temp_mem[1983];

   memory[496][0] = temp_mem[1984];
   memory[496][1] = temp_mem[1985];
   memory[496][2] = temp_mem[1986];
   memory[496][3] = temp_mem[1987];

   memory[497][0] = temp_mem[1988];
   memory[497][1] = temp_mem[1989];
   memory[497][2] = temp_mem[1990];
   memory[497][3] = temp_mem[1991];

   memory[498][0] = temp_mem[1992];
   memory[498][1] = temp_mem[1993];
   memory[498][2] = temp_mem[1994];
   memory[498][3] = temp_mem[1995];

   memory[499][0] = temp_mem[1996];
   memory[499][1] = temp_mem[1997];
   memory[499][2] = temp_mem[1998];
   memory[499][3] = temp_mem[1999];

   memory[500][0] = temp_mem[2000];
   memory[500][1] = temp_mem[2001];
   memory[500][2] = temp_mem[2002];
   memory[500][3] = temp_mem[2003];

   memory[501][0] = temp_mem[2004];
   memory[501][1] = temp_mem[2005];
   memory[501][2] = temp_mem[2006];
   memory[501][3] = temp_mem[2007];

   memory[502][0] = temp_mem[2008];
   memory[502][1] = temp_mem[2009];
   memory[502][2] = temp_mem[2010];
   memory[502][3] = temp_mem[2011];

   memory[503][0] = temp_mem[2012];
   memory[503][1] = temp_mem[2013];
   memory[503][2] = temp_mem[2014];
   memory[503][3] = temp_mem[2015];

   memory[504][0] = temp_mem[2016];
   memory[504][1] = temp_mem[2017];
   memory[504][2] = temp_mem[2018];
   memory[504][3] = temp_mem[2019];

   memory[505][0] = temp_mem[2020];
   memory[505][1] = temp_mem[2021];
   memory[505][2] = temp_mem[2022];
   memory[505][3] = temp_mem[2023];

   memory[506][0] = temp_mem[2024];
   memory[506][1] = temp_mem[2025];
   memory[506][2] = temp_mem[2026];
   memory[506][3] = temp_mem[2027];

   memory[507][0] = temp_mem[2028];
   memory[507][1] = temp_mem[2029];
   memory[507][2] = temp_mem[2030];
   memory[507][3] = temp_mem[2031];

   memory[508][0] = temp_mem[2032];
   memory[508][1] = temp_mem[2033];
   memory[508][2] = temp_mem[2034];
   memory[508][3] = temp_mem[2035];

   memory[509][0] = temp_mem[2036];
   memory[509][1] = temp_mem[2037];
   memory[509][2] = temp_mem[2038];
   memory[509][3] = temp_mem[2039];

   memory[510][0] = temp_mem[2040];
   memory[510][1] = temp_mem[2041];
   memory[510][2] = temp_mem[2042];
   memory[510][3] = temp_mem[2043];

   memory[511][0] = temp_mem[2044];
   memory[511][1] = temp_mem[2045];
   memory[511][2] = temp_mem[2046];
   memory[511][3] = temp_mem[2047];

   memory[512][0] = temp_mem[2048];
   memory[512][1] = temp_mem[2049];
   memory[512][2] = temp_mem[2050];
   memory[512][3] = temp_mem[2051];

   memory[513][0] = temp_mem[2052];
   memory[513][1] = temp_mem[2053];
   memory[513][2] = temp_mem[2054];
   memory[513][3] = temp_mem[2055];

   memory[514][0] = temp_mem[2056];
   memory[514][1] = temp_mem[2057];
   memory[514][2] = temp_mem[2058];
   memory[514][3] = temp_mem[2059];

   memory[515][0] = temp_mem[2060];
   memory[515][1] = temp_mem[2061];
   memory[515][2] = temp_mem[2062];
   memory[515][3] = temp_mem[2063];

   memory[516][0] = temp_mem[2064];
   memory[516][1] = temp_mem[2065];
   memory[516][2] = temp_mem[2066];
   memory[516][3] = temp_mem[2067];

   memory[517][0] = temp_mem[2068];
   memory[517][1] = temp_mem[2069];
   memory[517][2] = temp_mem[2070];
   memory[517][3] = temp_mem[2071];

   memory[518][0] = temp_mem[2072];
   memory[518][1] = temp_mem[2073];
   memory[518][2] = temp_mem[2074];
   memory[518][3] = temp_mem[2075];

   memory[519][0] = temp_mem[2076];
   memory[519][1] = temp_mem[2077];
   memory[519][2] = temp_mem[2078];
   memory[519][3] = temp_mem[2079];

   memory[520][0] = temp_mem[2080];
   memory[520][1] = temp_mem[2081];
   memory[520][2] = temp_mem[2082];
   memory[520][3] = temp_mem[2083];

   memory[521][0] = temp_mem[2084];
   memory[521][1] = temp_mem[2085];
   memory[521][2] = temp_mem[2086];
   memory[521][3] = temp_mem[2087];

   memory[522][0] = temp_mem[2088];
   memory[522][1] = temp_mem[2089];
   memory[522][2] = temp_mem[2090];
   memory[522][3] = temp_mem[2091];

   memory[523][0] = temp_mem[2092];
   memory[523][1] = temp_mem[2093];
   memory[523][2] = temp_mem[2094];
   memory[523][3] = temp_mem[2095];

   memory[524][0] = temp_mem[2096];
   memory[524][1] = temp_mem[2097];
   memory[524][2] = temp_mem[2098];
   memory[524][3] = temp_mem[2099];

   memory[525][0] = temp_mem[2100];
   memory[525][1] = temp_mem[2101];
   memory[525][2] = temp_mem[2102];
   memory[525][3] = temp_mem[2103];

   memory[526][0] = temp_mem[2104];
   memory[526][1] = temp_mem[2105];
   memory[526][2] = temp_mem[2106];
   memory[526][3] = temp_mem[2107];

   memory[527][0] = temp_mem[2108];
   memory[527][1] = temp_mem[2109];
   memory[527][2] = temp_mem[2110];
   memory[527][3] = temp_mem[2111];

   memory[528][0] = temp_mem[2112];
   memory[528][1] = temp_mem[2113];
   memory[528][2] = temp_mem[2114];
   memory[528][3] = temp_mem[2115];

   memory[529][0] = temp_mem[2116];
   memory[529][1] = temp_mem[2117];
   memory[529][2] = temp_mem[2118];
   memory[529][3] = temp_mem[2119];

   memory[530][0] = temp_mem[2120];
   memory[530][1] = temp_mem[2121];
   memory[530][2] = temp_mem[2122];
   memory[530][3] = temp_mem[2123];

   memory[531][0] = temp_mem[2124];
   memory[531][1] = temp_mem[2125];
   memory[531][2] = temp_mem[2126];
   memory[531][3] = temp_mem[2127];

   memory[532][0] = temp_mem[2128];
   memory[532][1] = temp_mem[2129];
   memory[532][2] = temp_mem[2130];
   memory[532][3] = temp_mem[2131];

   memory[533][0] = temp_mem[2132];
   memory[533][1] = temp_mem[2133];
   memory[533][2] = temp_mem[2134];
   memory[533][3] = temp_mem[2135];

   memory[534][0] = temp_mem[2136];
   memory[534][1] = temp_mem[2137];
   memory[534][2] = temp_mem[2138];
   memory[534][3] = temp_mem[2139];

   memory[535][0] = temp_mem[2140];
   memory[535][1] = temp_mem[2141];
   memory[535][2] = temp_mem[2142];
   memory[535][3] = temp_mem[2143];

   memory[536][0] = temp_mem[2144];
   memory[536][1] = temp_mem[2145];
   memory[536][2] = temp_mem[2146];
   memory[536][3] = temp_mem[2147];

   memory[537][0] = temp_mem[2148];
   memory[537][1] = temp_mem[2149];
   memory[537][2] = temp_mem[2150];
   memory[537][3] = temp_mem[2151];

   memory[538][0] = temp_mem[2152];
   memory[538][1] = temp_mem[2153];
   memory[538][2] = temp_mem[2154];
   memory[538][3] = temp_mem[2155];

   memory[539][0] = temp_mem[2156];
   memory[539][1] = temp_mem[2157];
   memory[539][2] = temp_mem[2158];
   memory[539][3] = temp_mem[2159];

   memory[540][0] = temp_mem[2160];
   memory[540][1] = temp_mem[2161];
   memory[540][2] = temp_mem[2162];
   memory[540][3] = temp_mem[2163];

   memory[541][0] = temp_mem[2164];
   memory[541][1] = temp_mem[2165];
   memory[541][2] = temp_mem[2166];
   memory[541][3] = temp_mem[2167];

   memory[542][0] = temp_mem[2168];
   memory[542][1] = temp_mem[2169];
   memory[542][2] = temp_mem[2170];
   memory[542][3] = temp_mem[2171];

   memory[543][0] = temp_mem[2172];
   memory[543][1] = temp_mem[2173];
   memory[543][2] = temp_mem[2174];
   memory[543][3] = temp_mem[2175];

   memory[544][0] = temp_mem[2176];
   memory[544][1] = temp_mem[2177];
   memory[544][2] = temp_mem[2178];
   memory[544][3] = temp_mem[2179];

   memory[545][0] = temp_mem[2180];
   memory[545][1] = temp_mem[2181];
   memory[545][2] = temp_mem[2182];
   memory[545][3] = temp_mem[2183];

   memory[546][0] = temp_mem[2184];
   memory[546][1] = temp_mem[2185];
   memory[546][2] = temp_mem[2186];
   memory[546][3] = temp_mem[2187];

   memory[547][0] = temp_mem[2188];
   memory[547][1] = temp_mem[2189];
   memory[547][2] = temp_mem[2190];
   memory[547][3] = temp_mem[2191];

   memory[548][0] = temp_mem[2192];
   memory[548][1] = temp_mem[2193];
   memory[548][2] = temp_mem[2194];
   memory[548][3] = temp_mem[2195];

   memory[549][0] = temp_mem[2196];
   memory[549][1] = temp_mem[2197];
   memory[549][2] = temp_mem[2198];
   memory[549][3] = temp_mem[2199];

   memory[550][0] = temp_mem[2200];
   memory[550][1] = temp_mem[2201];
   memory[550][2] = temp_mem[2202];
   memory[550][3] = temp_mem[2203];

   memory[551][0] = temp_mem[2204];
   memory[551][1] = temp_mem[2205];
   memory[551][2] = temp_mem[2206];
   memory[551][3] = temp_mem[2207];

   memory[552][0] = temp_mem[2208];
   memory[552][1] = temp_mem[2209];
   memory[552][2] = temp_mem[2210];
   memory[552][3] = temp_mem[2211];

   memory[553][0] = temp_mem[2212];
   memory[553][1] = temp_mem[2213];
   memory[553][2] = temp_mem[2214];
   memory[553][3] = temp_mem[2215];

   memory[554][0] = temp_mem[2216];
   memory[554][1] = temp_mem[2217];
   memory[554][2] = temp_mem[2218];
   memory[554][3] = temp_mem[2219];

   memory[555][0] = temp_mem[2220];
   memory[555][1] = temp_mem[2221];
   memory[555][2] = temp_mem[2222];
   memory[555][3] = temp_mem[2223];

   memory[556][0] = temp_mem[2224];
   memory[556][1] = temp_mem[2225];
   memory[556][2] = temp_mem[2226];
   memory[556][3] = temp_mem[2227];

   memory[557][0] = temp_mem[2228];
   memory[557][1] = temp_mem[2229];
   memory[557][2] = temp_mem[2230];
   memory[557][3] = temp_mem[2231];

   memory[558][0] = temp_mem[2232];
   memory[558][1] = temp_mem[2233];
   memory[558][2] = temp_mem[2234];
   memory[558][3] = temp_mem[2235];

   memory[559][0] = temp_mem[2236];
   memory[559][1] = temp_mem[2237];
   memory[559][2] = temp_mem[2238];
   memory[559][3] = temp_mem[2239];

   memory[560][0] = temp_mem[2240];
   memory[560][1] = temp_mem[2241];
   memory[560][2] = temp_mem[2242];
   memory[560][3] = temp_mem[2243];

   memory[561][0] = temp_mem[2244];
   memory[561][1] = temp_mem[2245];
   memory[561][2] = temp_mem[2246];
   memory[561][3] = temp_mem[2247];

   memory[562][0] = temp_mem[2248];
   memory[562][1] = temp_mem[2249];
   memory[562][2] = temp_mem[2250];
   memory[562][3] = temp_mem[2251];

   memory[563][0] = temp_mem[2252];
   memory[563][1] = temp_mem[2253];
   memory[563][2] = temp_mem[2254];
   memory[563][3] = temp_mem[2255];

   memory[564][0] = temp_mem[2256];
   memory[564][1] = temp_mem[2257];
   memory[564][2] = temp_mem[2258];
   memory[564][3] = temp_mem[2259];

   memory[565][0] = temp_mem[2260];
   memory[565][1] = temp_mem[2261];
   memory[565][2] = temp_mem[2262];
   memory[565][3] = temp_mem[2263];

   memory[566][0] = temp_mem[2264];
   memory[566][1] = temp_mem[2265];
   memory[566][2] = temp_mem[2266];
   memory[566][3] = temp_mem[2267];

   memory[567][0] = temp_mem[2268];
   memory[567][1] = temp_mem[2269];
   memory[567][2] = temp_mem[2270];
   memory[567][3] = temp_mem[2271];

   memory[568][0] = temp_mem[2272];
   memory[568][1] = temp_mem[2273];
   memory[568][2] = temp_mem[2274];
   memory[568][3] = temp_mem[2275];

   memory[569][0] = temp_mem[2276];
   memory[569][1] = temp_mem[2277];
   memory[569][2] = temp_mem[2278];
   memory[569][3] = temp_mem[2279];

   memory[570][0] = temp_mem[2280];
   memory[570][1] = temp_mem[2281];
   memory[570][2] = temp_mem[2282];
   memory[570][3] = temp_mem[2283];

   memory[571][0] = temp_mem[2284];
   memory[571][1] = temp_mem[2285];
   memory[571][2] = temp_mem[2286];
   memory[571][3] = temp_mem[2287];

   memory[572][0] = temp_mem[2288];
   memory[572][1] = temp_mem[2289];
   memory[572][2] = temp_mem[2290];
   memory[572][3] = temp_mem[2291];

   memory[573][0] = temp_mem[2292];
   memory[573][1] = temp_mem[2293];
   memory[573][2] = temp_mem[2294];
   memory[573][3] = temp_mem[2295];

   memory[574][0] = temp_mem[2296];
   memory[574][1] = temp_mem[2297];
   memory[574][2] = temp_mem[2298];
   memory[574][3] = temp_mem[2299];

   memory[575][0] = temp_mem[2300];
   memory[575][1] = temp_mem[2301];
   memory[575][2] = temp_mem[2302];
   memory[575][3] = temp_mem[2303];

   memory[576][0] = temp_mem[2304];
   memory[576][1] = temp_mem[2305];
   memory[576][2] = temp_mem[2306];
   memory[576][3] = temp_mem[2307];

   memory[577][0] = temp_mem[2308];
   memory[577][1] = temp_mem[2309];
   memory[577][2] = temp_mem[2310];
   memory[577][3] = temp_mem[2311];

   memory[578][0] = temp_mem[2312];
   memory[578][1] = temp_mem[2313];
   memory[578][2] = temp_mem[2314];
   memory[578][3] = temp_mem[2315];

   memory[579][0] = temp_mem[2316];
   memory[579][1] = temp_mem[2317];
   memory[579][2] = temp_mem[2318];
   memory[579][3] = temp_mem[2319];

   memory[580][0] = temp_mem[2320];
   memory[580][1] = temp_mem[2321];
   memory[580][2] = temp_mem[2322];
   memory[580][3] = temp_mem[2323];

   memory[581][0] = temp_mem[2324];
   memory[581][1] = temp_mem[2325];
   memory[581][2] = temp_mem[2326];
   memory[581][3] = temp_mem[2327];

   memory[582][0] = temp_mem[2328];
   memory[582][1] = temp_mem[2329];
   memory[582][2] = temp_mem[2330];
   memory[582][3] = temp_mem[2331];

   memory[583][0] = temp_mem[2332];
   memory[583][1] = temp_mem[2333];
   memory[583][2] = temp_mem[2334];
   memory[583][3] = temp_mem[2335];

   memory[584][0] = temp_mem[2336];
   memory[584][1] = temp_mem[2337];
   memory[584][2] = temp_mem[2338];
   memory[584][3] = temp_mem[2339];

   memory[585][0] = temp_mem[2340];
   memory[585][1] = temp_mem[2341];
   memory[585][2] = temp_mem[2342];
   memory[585][3] = temp_mem[2343];

   memory[586][0] = temp_mem[2344];
   memory[586][1] = temp_mem[2345];
   memory[586][2] = temp_mem[2346];
   memory[586][3] = temp_mem[2347];

   memory[587][0] = temp_mem[2348];
   memory[587][1] = temp_mem[2349];
   memory[587][2] = temp_mem[2350];
   memory[587][3] = temp_mem[2351];

   memory[588][0] = temp_mem[2352];
   memory[588][1] = temp_mem[2353];
   memory[588][2] = temp_mem[2354];
   memory[588][3] = temp_mem[2355];

   memory[589][0] = temp_mem[2356];
   memory[589][1] = temp_mem[2357];
   memory[589][2] = temp_mem[2358];
   memory[589][3] = temp_mem[2359];

   memory[590][0] = temp_mem[2360];
   memory[590][1] = temp_mem[2361];
   memory[590][2] = temp_mem[2362];
   memory[590][3] = temp_mem[2363];

   memory[591][0] = temp_mem[2364];
   memory[591][1] = temp_mem[2365];
   memory[591][2] = temp_mem[2366];
   memory[591][3] = temp_mem[2367];

   memory[592][0] = temp_mem[2368];
   memory[592][1] = temp_mem[2369];
   memory[592][2] = temp_mem[2370];
   memory[592][3] = temp_mem[2371];

   memory[593][0] = temp_mem[2372];
   memory[593][1] = temp_mem[2373];
   memory[593][2] = temp_mem[2374];
   memory[593][3] = temp_mem[2375];

   memory[594][0] = temp_mem[2376];
   memory[594][1] = temp_mem[2377];
   memory[594][2] = temp_mem[2378];
   memory[594][3] = temp_mem[2379];

   memory[595][0] = temp_mem[2380];
   memory[595][1] = temp_mem[2381];
   memory[595][2] = temp_mem[2382];
   memory[595][3] = temp_mem[2383];

   memory[596][0] = temp_mem[2384];
   memory[596][1] = temp_mem[2385];
   memory[596][2] = temp_mem[2386];
   memory[596][3] = temp_mem[2387];

   memory[597][0] = temp_mem[2388];
   memory[597][1] = temp_mem[2389];
   memory[597][2] = temp_mem[2390];
   memory[597][3] = temp_mem[2391];

   memory[598][0] = temp_mem[2392];
   memory[598][1] = temp_mem[2393];
   memory[598][2] = temp_mem[2394];
   memory[598][3] = temp_mem[2395];

   memory[599][0] = temp_mem[2396];
   memory[599][1] = temp_mem[2397];
   memory[599][2] = temp_mem[2398];
   memory[599][3] = temp_mem[2399];

   memory[600][0] = temp_mem[2400];
   memory[600][1] = temp_mem[2401];
   memory[600][2] = temp_mem[2402];
   memory[600][3] = temp_mem[2403];

   memory[601][0] = temp_mem[2404];
   memory[601][1] = temp_mem[2405];
   memory[601][2] = temp_mem[2406];
   memory[601][3] = temp_mem[2407];

   memory[602][0] = temp_mem[2408];
   memory[602][1] = temp_mem[2409];
   memory[602][2] = temp_mem[2410];
   memory[602][3] = temp_mem[2411];

   memory[603][0] = temp_mem[2412];
   memory[603][1] = temp_mem[2413];
   memory[603][2] = temp_mem[2414];
   memory[603][3] = temp_mem[2415];

   memory[604][0] = temp_mem[2416];
   memory[604][1] = temp_mem[2417];
   memory[604][2] = temp_mem[2418];
   memory[604][3] = temp_mem[2419];

   memory[605][0] = temp_mem[2420];
   memory[605][1] = temp_mem[2421];
   memory[605][2] = temp_mem[2422];
   memory[605][3] = temp_mem[2423];

   memory[606][0] = temp_mem[2424];
   memory[606][1] = temp_mem[2425];
   memory[606][2] = temp_mem[2426];
   memory[606][3] = temp_mem[2427];

   memory[607][0] = temp_mem[2428];
   memory[607][1] = temp_mem[2429];
   memory[607][2] = temp_mem[2430];
   memory[607][3] = temp_mem[2431];

   memory[608][0] = temp_mem[2432];
   memory[608][1] = temp_mem[2433];
   memory[608][2] = temp_mem[2434];
   memory[608][3] = temp_mem[2435];

   memory[609][0] = temp_mem[2436];
   memory[609][1] = temp_mem[2437];
   memory[609][2] = temp_mem[2438];
   memory[609][3] = temp_mem[2439];

   memory[610][0] = temp_mem[2440];
   memory[610][1] = temp_mem[2441];
   memory[610][2] = temp_mem[2442];
   memory[610][3] = temp_mem[2443];

   memory[611][0] = temp_mem[2444];
   memory[611][1] = temp_mem[2445];
   memory[611][2] = temp_mem[2446];
   memory[611][3] = temp_mem[2447];

   memory[612][0] = temp_mem[2448];
   memory[612][1] = temp_mem[2449];
   memory[612][2] = temp_mem[2450];
   memory[612][3] = temp_mem[2451];

   memory[613][0] = temp_mem[2452];
   memory[613][1] = temp_mem[2453];
   memory[613][2] = temp_mem[2454];
   memory[613][3] = temp_mem[2455];

   memory[614][0] = temp_mem[2456];
   memory[614][1] = temp_mem[2457];
   memory[614][2] = temp_mem[2458];
   memory[614][3] = temp_mem[2459];

   memory[615][0] = temp_mem[2460];
   memory[615][1] = temp_mem[2461];
   memory[615][2] = temp_mem[2462];
   memory[615][3] = temp_mem[2463];

   memory[616][0] = temp_mem[2464];
   memory[616][1] = temp_mem[2465];
   memory[616][2] = temp_mem[2466];
   memory[616][3] = temp_mem[2467];

   memory[617][0] = temp_mem[2468];
   memory[617][1] = temp_mem[2469];
   memory[617][2] = temp_mem[2470];
   memory[617][3] = temp_mem[2471];

   memory[618][0] = temp_mem[2472];
   memory[618][1] = temp_mem[2473];
   memory[618][2] = temp_mem[2474];
   memory[618][3] = temp_mem[2475];

   memory[619][0] = temp_mem[2476];
   memory[619][1] = temp_mem[2477];
   memory[619][2] = temp_mem[2478];
   memory[619][3] = temp_mem[2479];

   memory[620][0] = temp_mem[2480];
   memory[620][1] = temp_mem[2481];
   memory[620][2] = temp_mem[2482];
   memory[620][3] = temp_mem[2483];

   memory[621][0] = temp_mem[2484];
   memory[621][1] = temp_mem[2485];
   memory[621][2] = temp_mem[2486];
   memory[621][3] = temp_mem[2487];

   memory[622][0] = temp_mem[2488];
   memory[622][1] = temp_mem[2489];
   memory[622][2] = temp_mem[2490];
   memory[622][3] = temp_mem[2491];

   memory[623][0] = temp_mem[2492];
   memory[623][1] = temp_mem[2493];
   memory[623][2] = temp_mem[2494];
   memory[623][3] = temp_mem[2495];

   memory[624][0] = temp_mem[2496];
   memory[624][1] = temp_mem[2497];
   memory[624][2] = temp_mem[2498];
   memory[624][3] = temp_mem[2499];

   memory[625][0] = temp_mem[2500];
   memory[625][1] = temp_mem[2501];
   memory[625][2] = temp_mem[2502];
   memory[625][3] = temp_mem[2503];

   memory[626][0] = temp_mem[2504];
   memory[626][1] = temp_mem[2505];
   memory[626][2] = temp_mem[2506];
   memory[626][3] = temp_mem[2507];

   memory[627][0] = temp_mem[2508];
   memory[627][1] = temp_mem[2509];
   memory[627][2] = temp_mem[2510];
   memory[627][3] = temp_mem[2511];

   memory[628][0] = temp_mem[2512];
   memory[628][1] = temp_mem[2513];
   memory[628][2] = temp_mem[2514];
   memory[628][3] = temp_mem[2515];

   memory[629][0] = temp_mem[2516];
   memory[629][1] = temp_mem[2517];
   memory[629][2] = temp_mem[2518];
   memory[629][3] = temp_mem[2519];

   memory[630][0] = temp_mem[2520];
   memory[630][1] = temp_mem[2521];
   memory[630][2] = temp_mem[2522];
   memory[630][3] = temp_mem[2523];

   memory[631][0] = temp_mem[2524];
   memory[631][1] = temp_mem[2525];
   memory[631][2] = temp_mem[2526];
   memory[631][3] = temp_mem[2527];

   memory[632][0] = temp_mem[2528];
   memory[632][1] = temp_mem[2529];
   memory[632][2] = temp_mem[2530];
   memory[632][3] = temp_mem[2531];

   memory[633][0] = temp_mem[2532];
   memory[633][1] = temp_mem[2533];
   memory[633][2] = temp_mem[2534];
   memory[633][3] = temp_mem[2535];

   memory[634][0] = temp_mem[2536];
   memory[634][1] = temp_mem[2537];
   memory[634][2] = temp_mem[2538];
   memory[634][3] = temp_mem[2539];

   memory[635][0] = temp_mem[2540];
   memory[635][1] = temp_mem[2541];
   memory[635][2] = temp_mem[2542];
   memory[635][3] = temp_mem[2543];

   memory[636][0] = temp_mem[2544];
   memory[636][1] = temp_mem[2545];
   memory[636][2] = temp_mem[2546];
   memory[636][3] = temp_mem[2547];

   memory[637][0] = temp_mem[2548];
   memory[637][1] = temp_mem[2549];
   memory[637][2] = temp_mem[2550];
   memory[637][3] = temp_mem[2551];

   memory[638][0] = temp_mem[2552];
   memory[638][1] = temp_mem[2553];
   memory[638][2] = temp_mem[2554];
   memory[638][3] = temp_mem[2555];

   memory[639][0] = temp_mem[2556];
   memory[639][1] = temp_mem[2557];
   memory[639][2] = temp_mem[2558];
   memory[639][3] = temp_mem[2559];

   memory[640][0] = temp_mem[2560];
   memory[640][1] = temp_mem[2561];
   memory[640][2] = temp_mem[2562];
   memory[640][3] = temp_mem[2563];

   memory[641][0] = temp_mem[2564];
   memory[641][1] = temp_mem[2565];
   memory[641][2] = temp_mem[2566];
   memory[641][3] = temp_mem[2567];

   memory[642][0] = temp_mem[2568];
   memory[642][1] = temp_mem[2569];
   memory[642][2] = temp_mem[2570];
   memory[642][3] = temp_mem[2571];

   memory[643][0] = temp_mem[2572];
   memory[643][1] = temp_mem[2573];
   memory[643][2] = temp_mem[2574];
   memory[643][3] = temp_mem[2575];

   memory[644][0] = temp_mem[2576];
   memory[644][1] = temp_mem[2577];
   memory[644][2] = temp_mem[2578];
   memory[644][3] = temp_mem[2579];

   memory[645][0] = temp_mem[2580];
   memory[645][1] = temp_mem[2581];
   memory[645][2] = temp_mem[2582];
   memory[645][3] = temp_mem[2583];

   memory[646][0] = temp_mem[2584];
   memory[646][1] = temp_mem[2585];
   memory[646][2] = temp_mem[2586];
   memory[646][3] = temp_mem[2587];

   memory[647][0] = temp_mem[2588];
   memory[647][1] = temp_mem[2589];
   memory[647][2] = temp_mem[2590];
   memory[647][3] = temp_mem[2591];

   memory[648][0] = temp_mem[2592];
   memory[648][1] = temp_mem[2593];
   memory[648][2] = temp_mem[2594];
   memory[648][3] = temp_mem[2595];

   memory[649][0] = temp_mem[2596];
   memory[649][1] = temp_mem[2597];
   memory[649][2] = temp_mem[2598];
   memory[649][3] = temp_mem[2599];

   memory[650][0] = temp_mem[2600];
   memory[650][1] = temp_mem[2601];
   memory[650][2] = temp_mem[2602];
   memory[650][3] = temp_mem[2603];

   memory[651][0] = temp_mem[2604];
   memory[651][1] = temp_mem[2605];
   memory[651][2] = temp_mem[2606];
   memory[651][3] = temp_mem[2607];

   memory[652][0] = temp_mem[2608];
   memory[652][1] = temp_mem[2609];
   memory[652][2] = temp_mem[2610];
   memory[652][3] = temp_mem[2611];

   memory[653][0] = temp_mem[2612];
   memory[653][1] = temp_mem[2613];
   memory[653][2] = temp_mem[2614];
   memory[653][3] = temp_mem[2615];

   memory[654][0] = temp_mem[2616];
   memory[654][1] = temp_mem[2617];
   memory[654][2] = temp_mem[2618];
   memory[654][3] = temp_mem[2619];

   memory[655][0] = temp_mem[2620];
   memory[655][1] = temp_mem[2621];
   memory[655][2] = temp_mem[2622];
   memory[655][3] = temp_mem[2623];

   memory[656][0] = temp_mem[2624];
   memory[656][1] = temp_mem[2625];
   memory[656][2] = temp_mem[2626];
   memory[656][3] = temp_mem[2627];

   memory[657][0] = temp_mem[2628];
   memory[657][1] = temp_mem[2629];
   memory[657][2] = temp_mem[2630];
   memory[657][3] = temp_mem[2631];

   memory[658][0] = temp_mem[2632];
   memory[658][1] = temp_mem[2633];
   memory[658][2] = temp_mem[2634];
   memory[658][3] = temp_mem[2635];

   memory[659][0] = temp_mem[2636];
   memory[659][1] = temp_mem[2637];
   memory[659][2] = temp_mem[2638];
   memory[659][3] = temp_mem[2639];

   memory[660][0] = temp_mem[2640];
   memory[660][1] = temp_mem[2641];
   memory[660][2] = temp_mem[2642];
   memory[660][3] = temp_mem[2643];

   memory[661][0] = temp_mem[2644];
   memory[661][1] = temp_mem[2645];
   memory[661][2] = temp_mem[2646];
   memory[661][3] = temp_mem[2647];

   memory[662][0] = temp_mem[2648];
   memory[662][1] = temp_mem[2649];
   memory[662][2] = temp_mem[2650];
   memory[662][3] = temp_mem[2651];

   memory[663][0] = temp_mem[2652];
   memory[663][1] = temp_mem[2653];
   memory[663][2] = temp_mem[2654];
   memory[663][3] = temp_mem[2655];

   memory[664][0] = temp_mem[2656];
   memory[664][1] = temp_mem[2657];
   memory[664][2] = temp_mem[2658];
   memory[664][3] = temp_mem[2659];

   memory[665][0] = temp_mem[2660];
   memory[665][1] = temp_mem[2661];
   memory[665][2] = temp_mem[2662];
   memory[665][3] = temp_mem[2663];

   memory[666][0] = temp_mem[2664];
   memory[666][1] = temp_mem[2665];
   memory[666][2] = temp_mem[2666];
   memory[666][3] = temp_mem[2667];

   memory[667][0] = temp_mem[2668];
   memory[667][1] = temp_mem[2669];
   memory[667][2] = temp_mem[2670];
   memory[667][3] = temp_mem[2671];

   memory[668][0] = temp_mem[2672];
   memory[668][1] = temp_mem[2673];
   memory[668][2] = temp_mem[2674];
   memory[668][3] = temp_mem[2675];

   memory[669][0] = temp_mem[2676];
   memory[669][1] = temp_mem[2677];
   memory[669][2] = temp_mem[2678];
   memory[669][3] = temp_mem[2679];

   memory[670][0] = temp_mem[2680];
   memory[670][1] = temp_mem[2681];
   memory[670][2] = temp_mem[2682];
   memory[670][3] = temp_mem[2683];

   memory[671][0] = temp_mem[2684];
   memory[671][1] = temp_mem[2685];
   memory[671][2] = temp_mem[2686];
   memory[671][3] = temp_mem[2687];

   memory[672][0] = temp_mem[2688];
   memory[672][1] = temp_mem[2689];
   memory[672][2] = temp_mem[2690];
   memory[672][3] = temp_mem[2691];

   memory[673][0] = temp_mem[2692];
   memory[673][1] = temp_mem[2693];
   memory[673][2] = temp_mem[2694];
   memory[673][3] = temp_mem[2695];

   memory[674][0] = temp_mem[2696];
   memory[674][1] = temp_mem[2697];
   memory[674][2] = temp_mem[2698];
   memory[674][3] = temp_mem[2699];

   memory[675][0] = temp_mem[2700];
   memory[675][1] = temp_mem[2701];
   memory[675][2] = temp_mem[2702];
   memory[675][3] = temp_mem[2703];

   memory[676][0] = temp_mem[2704];
   memory[676][1] = temp_mem[2705];
   memory[676][2] = temp_mem[2706];
   memory[676][3] = temp_mem[2707];

   memory[677][0] = temp_mem[2708];
   memory[677][1] = temp_mem[2709];
   memory[677][2] = temp_mem[2710];
   memory[677][3] = temp_mem[2711];

   memory[678][0] = temp_mem[2712];
   memory[678][1] = temp_mem[2713];
   memory[678][2] = temp_mem[2714];
   memory[678][3] = temp_mem[2715];

   memory[679][0] = temp_mem[2716];
   memory[679][1] = temp_mem[2717];
   memory[679][2] = temp_mem[2718];
   memory[679][3] = temp_mem[2719];

   memory[680][0] = temp_mem[2720];
   memory[680][1] = temp_mem[2721];
   memory[680][2] = temp_mem[2722];
   memory[680][3] = temp_mem[2723];

   memory[681][0] = temp_mem[2724];
   memory[681][1] = temp_mem[2725];
   memory[681][2] = temp_mem[2726];
   memory[681][3] = temp_mem[2727];

   memory[682][0] = temp_mem[2728];
   memory[682][1] = temp_mem[2729];
   memory[682][2] = temp_mem[2730];
   memory[682][3] = temp_mem[2731];

   memory[683][0] = temp_mem[2732];
   memory[683][1] = temp_mem[2733];
   memory[683][2] = temp_mem[2734];
   memory[683][3] = temp_mem[2735];

   memory[684][0] = temp_mem[2736];
   memory[684][1] = temp_mem[2737];
   memory[684][2] = temp_mem[2738];
   memory[684][3] = temp_mem[2739];

   memory[685][0] = temp_mem[2740];
   memory[685][1] = temp_mem[2741];
   memory[685][2] = temp_mem[2742];
   memory[685][3] = temp_mem[2743];

   memory[686][0] = temp_mem[2744];
   memory[686][1] = temp_mem[2745];
   memory[686][2] = temp_mem[2746];
   memory[686][3] = temp_mem[2747];

   memory[687][0] = temp_mem[2748];
   memory[687][1] = temp_mem[2749];
   memory[687][2] = temp_mem[2750];
   memory[687][3] = temp_mem[2751];

   memory[688][0] = temp_mem[2752];
   memory[688][1] = temp_mem[2753];
   memory[688][2] = temp_mem[2754];
   memory[688][3] = temp_mem[2755];

   memory[689][0] = temp_mem[2756];
   memory[689][1] = temp_mem[2757];
   memory[689][2] = temp_mem[2758];
   memory[689][3] = temp_mem[2759];

   memory[690][0] = temp_mem[2760];
   memory[690][1] = temp_mem[2761];
   memory[690][2] = temp_mem[2762];
   memory[690][3] = temp_mem[2763];

   memory[691][0] = temp_mem[2764];
   memory[691][1] = temp_mem[2765];
   memory[691][2] = temp_mem[2766];
   memory[691][3] = temp_mem[2767];

   memory[692][0] = temp_mem[2768];
   memory[692][1] = temp_mem[2769];
   memory[692][2] = temp_mem[2770];
   memory[692][3] = temp_mem[2771];

   memory[693][0] = temp_mem[2772];
   memory[693][1] = temp_mem[2773];
   memory[693][2] = temp_mem[2774];
   memory[693][3] = temp_mem[2775];

   memory[694][0] = temp_mem[2776];
   memory[694][1] = temp_mem[2777];
   memory[694][2] = temp_mem[2778];
   memory[694][3] = temp_mem[2779];

   memory[695][0] = temp_mem[2780];
   memory[695][1] = temp_mem[2781];
   memory[695][2] = temp_mem[2782];
   memory[695][3] = temp_mem[2783];

   memory[696][0] = temp_mem[2784];
   memory[696][1] = temp_mem[2785];
   memory[696][2] = temp_mem[2786];
   memory[696][3] = temp_mem[2787];

   memory[697][0] = temp_mem[2788];
   memory[697][1] = temp_mem[2789];
   memory[697][2] = temp_mem[2790];
   memory[697][3] = temp_mem[2791];

   memory[698][0] = temp_mem[2792];
   memory[698][1] = temp_mem[2793];
   memory[698][2] = temp_mem[2794];
   memory[698][3] = temp_mem[2795];

   memory[699][0] = temp_mem[2796];
   memory[699][1] = temp_mem[2797];
   memory[699][2] = temp_mem[2798];
   memory[699][3] = temp_mem[2799];

   memory[700][0] = temp_mem[2800];
   memory[700][1] = temp_mem[2801];
   memory[700][2] = temp_mem[2802];
   memory[700][3] = temp_mem[2803];

   memory[701][0] = temp_mem[2804];
   memory[701][1] = temp_mem[2805];
   memory[701][2] = temp_mem[2806];
   memory[701][3] = temp_mem[2807];

   memory[702][0] = temp_mem[2808];
   memory[702][1] = temp_mem[2809];
   memory[702][2] = temp_mem[2810];
   memory[702][3] = temp_mem[2811];

   memory[703][0] = temp_mem[2812];
   memory[703][1] = temp_mem[2813];
   memory[703][2] = temp_mem[2814];
   memory[703][3] = temp_mem[2815];

   memory[704][0] = temp_mem[2816];
   memory[704][1] = temp_mem[2817];
   memory[704][2] = temp_mem[2818];
   memory[704][3] = temp_mem[2819];

   memory[705][0] = temp_mem[2820];
   memory[705][1] = temp_mem[2821];
   memory[705][2] = temp_mem[2822];
   memory[705][3] = temp_mem[2823];

   memory[706][0] = temp_mem[2824];
   memory[706][1] = temp_mem[2825];
   memory[706][2] = temp_mem[2826];
   memory[706][3] = temp_mem[2827];

   memory[707][0] = temp_mem[2828];
   memory[707][1] = temp_mem[2829];
   memory[707][2] = temp_mem[2830];
   memory[707][3] = temp_mem[2831];

   memory[708][0] = temp_mem[2832];
   memory[708][1] = temp_mem[2833];
   memory[708][2] = temp_mem[2834];
   memory[708][3] = temp_mem[2835];

   memory[709][0] = temp_mem[2836];
   memory[709][1] = temp_mem[2837];
   memory[709][2] = temp_mem[2838];
   memory[709][3] = temp_mem[2839];

   memory[710][0] = temp_mem[2840];
   memory[710][1] = temp_mem[2841];
   memory[710][2] = temp_mem[2842];
   memory[710][3] = temp_mem[2843];

   memory[711][0] = temp_mem[2844];
   memory[711][1] = temp_mem[2845];
   memory[711][2] = temp_mem[2846];
   memory[711][3] = temp_mem[2847];

   memory[712][0] = temp_mem[2848];
   memory[712][1] = temp_mem[2849];
   memory[712][2] = temp_mem[2850];
   memory[712][3] = temp_mem[2851];

   memory[713][0] = temp_mem[2852];
   memory[713][1] = temp_mem[2853];
   memory[713][2] = temp_mem[2854];
   memory[713][3] = temp_mem[2855];

   memory[714][0] = temp_mem[2856];
   memory[714][1] = temp_mem[2857];
   memory[714][2] = temp_mem[2858];
   memory[714][3] = temp_mem[2859];

   memory[715][0] = temp_mem[2860];
   memory[715][1] = temp_mem[2861];
   memory[715][2] = temp_mem[2862];
   memory[715][3] = temp_mem[2863];

   memory[716][0] = temp_mem[2864];
   memory[716][1] = temp_mem[2865];
   memory[716][2] = temp_mem[2866];
   memory[716][3] = temp_mem[2867];

   memory[717][0] = temp_mem[2868];
   memory[717][1] = temp_mem[2869];
   memory[717][2] = temp_mem[2870];
   memory[717][3] = temp_mem[2871];

   memory[718][0] = temp_mem[2872];
   memory[718][1] = temp_mem[2873];
   memory[718][2] = temp_mem[2874];
   memory[718][3] = temp_mem[2875];

   memory[719][0] = temp_mem[2876];
   memory[719][1] = temp_mem[2877];
   memory[719][2] = temp_mem[2878];
   memory[719][3] = temp_mem[2879];

   memory[720][0] = temp_mem[2880];
   memory[720][1] = temp_mem[2881];
   memory[720][2] = temp_mem[2882];
   memory[720][3] = temp_mem[2883];

   memory[721][0] = temp_mem[2884];
   memory[721][1] = temp_mem[2885];
   memory[721][2] = temp_mem[2886];
   memory[721][3] = temp_mem[2887];

   memory[722][0] = temp_mem[2888];
   memory[722][1] = temp_mem[2889];
   memory[722][2] = temp_mem[2890];
   memory[722][3] = temp_mem[2891];

   memory[723][0] = temp_mem[2892];
   memory[723][1] = temp_mem[2893];
   memory[723][2] = temp_mem[2894];
   memory[723][3] = temp_mem[2895];

   memory[724][0] = temp_mem[2896];
   memory[724][1] = temp_mem[2897];
   memory[724][2] = temp_mem[2898];
   memory[724][3] = temp_mem[2899];

   memory[725][0] = temp_mem[2900];
   memory[725][1] = temp_mem[2901];
   memory[725][2] = temp_mem[2902];
   memory[725][3] = temp_mem[2903];

   memory[726][0] = temp_mem[2904];
   memory[726][1] = temp_mem[2905];
   memory[726][2] = temp_mem[2906];
   memory[726][3] = temp_mem[2907];

   memory[727][0] = temp_mem[2908];
   memory[727][1] = temp_mem[2909];
   memory[727][2] = temp_mem[2910];
   memory[727][3] = temp_mem[2911];

   memory[728][0] = temp_mem[2912];
   memory[728][1] = temp_mem[2913];
   memory[728][2] = temp_mem[2914];
   memory[728][3] = temp_mem[2915];

   memory[729][0] = temp_mem[2916];
   memory[729][1] = temp_mem[2917];
   memory[729][2] = temp_mem[2918];
   memory[729][3] = temp_mem[2919];

   memory[730][0] = temp_mem[2920];
   memory[730][1] = temp_mem[2921];
   memory[730][2] = temp_mem[2922];
   memory[730][3] = temp_mem[2923];

   memory[731][0] = temp_mem[2924];
   memory[731][1] = temp_mem[2925];
   memory[731][2] = temp_mem[2926];
   memory[731][3] = temp_mem[2927];

   memory[732][0] = temp_mem[2928];
   memory[732][1] = temp_mem[2929];
   memory[732][2] = temp_mem[2930];
   memory[732][3] = temp_mem[2931];

   memory[733][0] = temp_mem[2932];
   memory[733][1] = temp_mem[2933];
   memory[733][2] = temp_mem[2934];
   memory[733][3] = temp_mem[2935];

   memory[734][0] = temp_mem[2936];
   memory[734][1] = temp_mem[2937];
   memory[734][2] = temp_mem[2938];
   memory[734][3] = temp_mem[2939];

   memory[735][0] = temp_mem[2940];
   memory[735][1] = temp_mem[2941];
   memory[735][2] = temp_mem[2942];
   memory[735][3] = temp_mem[2943];

   memory[736][0] = temp_mem[2944];
   memory[736][1] = temp_mem[2945];
   memory[736][2] = temp_mem[2946];
   memory[736][3] = temp_mem[2947];

   memory[737][0] = temp_mem[2948];
   memory[737][1] = temp_mem[2949];
   memory[737][2] = temp_mem[2950];
   memory[737][3] = temp_mem[2951];

   memory[738][0] = temp_mem[2952];
   memory[738][1] = temp_mem[2953];
   memory[738][2] = temp_mem[2954];
   memory[738][3] = temp_mem[2955];

   memory[739][0] = temp_mem[2956];
   memory[739][1] = temp_mem[2957];
   memory[739][2] = temp_mem[2958];
   memory[739][3] = temp_mem[2959];

   memory[740][0] = temp_mem[2960];
   memory[740][1] = temp_mem[2961];
   memory[740][2] = temp_mem[2962];
   memory[740][3] = temp_mem[2963];

   memory[741][0] = temp_mem[2964];
   memory[741][1] = temp_mem[2965];
   memory[741][2] = temp_mem[2966];
   memory[741][3] = temp_mem[2967];

   memory[742][0] = temp_mem[2968];
   memory[742][1] = temp_mem[2969];
   memory[742][2] = temp_mem[2970];
   memory[742][3] = temp_mem[2971];

   memory[743][0] = temp_mem[2972];
   memory[743][1] = temp_mem[2973];
   memory[743][2] = temp_mem[2974];
   memory[743][3] = temp_mem[2975];

   memory[744][0] = temp_mem[2976];
   memory[744][1] = temp_mem[2977];
   memory[744][2] = temp_mem[2978];
   memory[744][3] = temp_mem[2979];

   memory[745][0] = temp_mem[2980];
   memory[745][1] = temp_mem[2981];
   memory[745][2] = temp_mem[2982];
   memory[745][3] = temp_mem[2983];

   memory[746][0] = temp_mem[2984];
   memory[746][1] = temp_mem[2985];
   memory[746][2] = temp_mem[2986];
   memory[746][3] = temp_mem[2987];

   memory[747][0] = temp_mem[2988];
   memory[747][1] = temp_mem[2989];
   memory[747][2] = temp_mem[2990];
   memory[747][3] = temp_mem[2991];

   memory[748][0] = temp_mem[2992];
   memory[748][1] = temp_mem[2993];
   memory[748][2] = temp_mem[2994];
   memory[748][3] = temp_mem[2995];

   memory[749][0] = temp_mem[2996];
   memory[749][1] = temp_mem[2997];
   memory[749][2] = temp_mem[2998];
   memory[749][3] = temp_mem[2999];

   memory[750][0] = temp_mem[3000];
   memory[750][1] = temp_mem[3001];
   memory[750][2] = temp_mem[3002];
   memory[750][3] = temp_mem[3003];

   memory[751][0] = temp_mem[3004];
   memory[751][1] = temp_mem[3005];
   memory[751][2] = temp_mem[3006];
   memory[751][3] = temp_mem[3007];

   memory[752][0] = temp_mem[3008];
   memory[752][1] = temp_mem[3009];
   memory[752][2] = temp_mem[3010];
   memory[752][3] = temp_mem[3011];

   memory[753][0] = temp_mem[3012];
   memory[753][1] = temp_mem[3013];
   memory[753][2] = temp_mem[3014];
   memory[753][3] = temp_mem[3015];

   memory[754][0] = temp_mem[3016];
   memory[754][1] = temp_mem[3017];
   memory[754][2] = temp_mem[3018];
   memory[754][3] = temp_mem[3019];

   memory[755][0] = temp_mem[3020];
   memory[755][1] = temp_mem[3021];
   memory[755][2] = temp_mem[3022];
   memory[755][3] = temp_mem[3023];

   memory[756][0] = temp_mem[3024];
   memory[756][1] = temp_mem[3025];
   memory[756][2] = temp_mem[3026];
   memory[756][3] = temp_mem[3027];

   memory[757][0] = temp_mem[3028];
   memory[757][1] = temp_mem[3029];
   memory[757][2] = temp_mem[3030];
   memory[757][3] = temp_mem[3031];

   memory[758][0] = temp_mem[3032];
   memory[758][1] = temp_mem[3033];
   memory[758][2] = temp_mem[3034];
   memory[758][3] = temp_mem[3035];

   memory[759][0] = temp_mem[3036];
   memory[759][1] = temp_mem[3037];
   memory[759][2] = temp_mem[3038];
   memory[759][3] = temp_mem[3039];

   memory[760][0] = temp_mem[3040];
   memory[760][1] = temp_mem[3041];
   memory[760][2] = temp_mem[3042];
   memory[760][3] = temp_mem[3043];

   memory[761][0] = temp_mem[3044];
   memory[761][1] = temp_mem[3045];
   memory[761][2] = temp_mem[3046];
   memory[761][3] = temp_mem[3047];

   memory[762][0] = temp_mem[3048];
   memory[762][1] = temp_mem[3049];
   memory[762][2] = temp_mem[3050];
   memory[762][3] = temp_mem[3051];

   memory[763][0] = temp_mem[3052];
   memory[763][1] = temp_mem[3053];
   memory[763][2] = temp_mem[3054];
   memory[763][3] = temp_mem[3055];

   memory[764][0] = temp_mem[3056];
   memory[764][1] = temp_mem[3057];
   memory[764][2] = temp_mem[3058];
   memory[764][3] = temp_mem[3059];

   memory[765][0] = temp_mem[3060];
   memory[765][1] = temp_mem[3061];
   memory[765][2] = temp_mem[3062];
   memory[765][3] = temp_mem[3063];

   memory[766][0] = temp_mem[3064];
   memory[766][1] = temp_mem[3065];
   memory[766][2] = temp_mem[3066];
   memory[766][3] = temp_mem[3067];

   memory[767][0] = temp_mem[3068];
   memory[767][1] = temp_mem[3069];
   memory[767][2] = temp_mem[3070];
   memory[767][3] = temp_mem[3071];

   memory[768][0] = temp_mem[3072];
   memory[768][1] = temp_mem[3073];
   memory[768][2] = temp_mem[3074];
   memory[768][3] = temp_mem[3075];

   memory[769][0] = temp_mem[3076];
   memory[769][1] = temp_mem[3077];
   memory[769][2] = temp_mem[3078];
   memory[769][3] = temp_mem[3079];

   memory[770][0] = temp_mem[3080];
   memory[770][1] = temp_mem[3081];
   memory[770][2] = temp_mem[3082];
   memory[770][3] = temp_mem[3083];

   memory[771][0] = temp_mem[3084];
   memory[771][1] = temp_mem[3085];
   memory[771][2] = temp_mem[3086];
   memory[771][3] = temp_mem[3087];

   memory[772][0] = temp_mem[3088];
   memory[772][1] = temp_mem[3089];
   memory[772][2] = temp_mem[3090];
   memory[772][3] = temp_mem[3091];

   memory[773][0] = temp_mem[3092];
   memory[773][1] = temp_mem[3093];
   memory[773][2] = temp_mem[3094];
   memory[773][3] = temp_mem[3095];

   memory[774][0] = temp_mem[3096];
   memory[774][1] = temp_mem[3097];
   memory[774][2] = temp_mem[3098];
   memory[774][3] = temp_mem[3099];

   memory[775][0] = temp_mem[3100];
   memory[775][1] = temp_mem[3101];
   memory[775][2] = temp_mem[3102];
   memory[775][3] = temp_mem[3103];

   memory[776][0] = temp_mem[3104];
   memory[776][1] = temp_mem[3105];
   memory[776][2] = temp_mem[3106];
   memory[776][3] = temp_mem[3107];

   memory[777][0] = temp_mem[3108];
   memory[777][1] = temp_mem[3109];
   memory[777][2] = temp_mem[3110];
   memory[777][3] = temp_mem[3111];

   memory[778][0] = temp_mem[3112];
   memory[778][1] = temp_mem[3113];
   memory[778][2] = temp_mem[3114];
   memory[778][3] = temp_mem[3115];

   memory[779][0] = temp_mem[3116];
   memory[779][1] = temp_mem[3117];
   memory[779][2] = temp_mem[3118];
   memory[779][3] = temp_mem[3119];

   memory[780][0] = temp_mem[3120];
   memory[780][1] = temp_mem[3121];
   memory[780][2] = temp_mem[3122];
   memory[780][3] = temp_mem[3123];

   memory[781][0] = temp_mem[3124];
   memory[781][1] = temp_mem[3125];
   memory[781][2] = temp_mem[3126];
   memory[781][3] = temp_mem[3127];

   memory[782][0] = temp_mem[3128];
   memory[782][1] = temp_mem[3129];
   memory[782][2] = temp_mem[3130];
   memory[782][3] = temp_mem[3131];

   memory[783][0] = temp_mem[3132];
   memory[783][1] = temp_mem[3133];
   memory[783][2] = temp_mem[3134];
   memory[783][3] = temp_mem[3135];

   memory[784][0] = temp_mem[3136];
   memory[784][1] = temp_mem[3137];
   memory[784][2] = temp_mem[3138];
   memory[784][3] = temp_mem[3139];

   memory[785][0] = temp_mem[3140];
   memory[785][1] = temp_mem[3141];
   memory[785][2] = temp_mem[3142];
   memory[785][3] = temp_mem[3143];

   memory[786][0] = temp_mem[3144];
   memory[786][1] = temp_mem[3145];
   memory[786][2] = temp_mem[3146];
   memory[786][3] = temp_mem[3147];

   memory[787][0] = temp_mem[3148];
   memory[787][1] = temp_mem[3149];
   memory[787][2] = temp_mem[3150];
   memory[787][3] = temp_mem[3151];

   memory[788][0] = temp_mem[3152];
   memory[788][1] = temp_mem[3153];
   memory[788][2] = temp_mem[3154];
   memory[788][3] = temp_mem[3155];

   memory[789][0] = temp_mem[3156];
   memory[789][1] = temp_mem[3157];
   memory[789][2] = temp_mem[3158];
   memory[789][3] = temp_mem[3159];

   memory[790][0] = temp_mem[3160];
   memory[790][1] = temp_mem[3161];
   memory[790][2] = temp_mem[3162];
   memory[790][3] = temp_mem[3163];

   memory[791][0] = temp_mem[3164];
   memory[791][1] = temp_mem[3165];
   memory[791][2] = temp_mem[3166];
   memory[791][3] = temp_mem[3167];

   memory[792][0] = temp_mem[3168];
   memory[792][1] = temp_mem[3169];
   memory[792][2] = temp_mem[3170];
   memory[792][3] = temp_mem[3171];

   memory[793][0] = temp_mem[3172];
   memory[793][1] = temp_mem[3173];
   memory[793][2] = temp_mem[3174];
   memory[793][3] = temp_mem[3175];

   memory[794][0] = temp_mem[3176];
   memory[794][1] = temp_mem[3177];
   memory[794][2] = temp_mem[3178];
   memory[794][3] = temp_mem[3179];

   memory[795][0] = temp_mem[3180];
   memory[795][1] = temp_mem[3181];
   memory[795][2] = temp_mem[3182];
   memory[795][3] = temp_mem[3183];

   memory[796][0] = temp_mem[3184];
   memory[796][1] = temp_mem[3185];
   memory[796][2] = temp_mem[3186];
   memory[796][3] = temp_mem[3187];

   memory[797][0] = temp_mem[3188];
   memory[797][1] = temp_mem[3189];
   memory[797][2] = temp_mem[3190];
   memory[797][3] = temp_mem[3191];

   memory[798][0] = temp_mem[3192];
   memory[798][1] = temp_mem[3193];
   memory[798][2] = temp_mem[3194];
   memory[798][3] = temp_mem[3195];

   memory[799][0] = temp_mem[3196];
   memory[799][1] = temp_mem[3197];
   memory[799][2] = temp_mem[3198];
   memory[799][3] = temp_mem[3199];

   memory[800][0] = temp_mem[3200];
   memory[800][1] = temp_mem[3201];
   memory[800][2] = temp_mem[3202];
   memory[800][3] = temp_mem[3203];

   memory[801][0] = temp_mem[3204];
   memory[801][1] = temp_mem[3205];
   memory[801][2] = temp_mem[3206];
   memory[801][3] = temp_mem[3207];

   memory[802][0] = temp_mem[3208];
   memory[802][1] = temp_mem[3209];
   memory[802][2] = temp_mem[3210];
   memory[802][3] = temp_mem[3211];

   memory[803][0] = temp_mem[3212];
   memory[803][1] = temp_mem[3213];
   memory[803][2] = temp_mem[3214];
   memory[803][3] = temp_mem[3215];

   memory[804][0] = temp_mem[3216];
   memory[804][1] = temp_mem[3217];
   memory[804][2] = temp_mem[3218];
   memory[804][3] = temp_mem[3219];

   memory[805][0] = temp_mem[3220];
   memory[805][1] = temp_mem[3221];
   memory[805][2] = temp_mem[3222];
   memory[805][3] = temp_mem[3223];

   memory[806][0] = temp_mem[3224];
   memory[806][1] = temp_mem[3225];
   memory[806][2] = temp_mem[3226];
   memory[806][3] = temp_mem[3227];

   memory[807][0] = temp_mem[3228];
   memory[807][1] = temp_mem[3229];
   memory[807][2] = temp_mem[3230];
   memory[807][3] = temp_mem[3231];

   memory[808][0] = temp_mem[3232];
   memory[808][1] = temp_mem[3233];
   memory[808][2] = temp_mem[3234];
   memory[808][3] = temp_mem[3235];

   memory[809][0] = temp_mem[3236];
   memory[809][1] = temp_mem[3237];
   memory[809][2] = temp_mem[3238];
   memory[809][3] = temp_mem[3239];

   memory[810][0] = temp_mem[3240];
   memory[810][1] = temp_mem[3241];
   memory[810][2] = temp_mem[3242];
   memory[810][3] = temp_mem[3243];

   memory[811][0] = temp_mem[3244];
   memory[811][1] = temp_mem[3245];
   memory[811][2] = temp_mem[3246];
   memory[811][3] = temp_mem[3247];

   memory[812][0] = temp_mem[3248];
   memory[812][1] = temp_mem[3249];
   memory[812][2] = temp_mem[3250];
   memory[812][3] = temp_mem[3251];

   memory[813][0] = temp_mem[3252];
   memory[813][1] = temp_mem[3253];
   memory[813][2] = temp_mem[3254];
   memory[813][3] = temp_mem[3255];

   memory[814][0] = temp_mem[3256];
   memory[814][1] = temp_mem[3257];
   memory[814][2] = temp_mem[3258];
   memory[814][3] = temp_mem[3259];

   memory[815][0] = temp_mem[3260];
   memory[815][1] = temp_mem[3261];
   memory[815][2] = temp_mem[3262];
   memory[815][3] = temp_mem[3263];

   memory[816][0] = temp_mem[3264];
   memory[816][1] = temp_mem[3265];
   memory[816][2] = temp_mem[3266];
   memory[816][3] = temp_mem[3267];

   memory[817][0] = temp_mem[3268];
   memory[817][1] = temp_mem[3269];
   memory[817][2] = temp_mem[3270];
   memory[817][3] = temp_mem[3271];

   memory[818][0] = temp_mem[3272];
   memory[818][1] = temp_mem[3273];
   memory[818][2] = temp_mem[3274];
   memory[818][3] = temp_mem[3275];

   memory[819][0] = temp_mem[3276];
   memory[819][1] = temp_mem[3277];
   memory[819][2] = temp_mem[3278];
   memory[819][3] = temp_mem[3279];

   memory[820][0] = temp_mem[3280];
   memory[820][1] = temp_mem[3281];
   memory[820][2] = temp_mem[3282];
   memory[820][3] = temp_mem[3283];

   memory[821][0] = temp_mem[3284];
   memory[821][1] = temp_mem[3285];
   memory[821][2] = temp_mem[3286];
   memory[821][3] = temp_mem[3287];

   memory[822][0] = temp_mem[3288];
   memory[822][1] = temp_mem[3289];
   memory[822][2] = temp_mem[3290];
   memory[822][3] = temp_mem[3291];

   memory[823][0] = temp_mem[3292];
   memory[823][1] = temp_mem[3293];
   memory[823][2] = temp_mem[3294];
   memory[823][3] = temp_mem[3295];

   memory[824][0] = temp_mem[3296];
   memory[824][1] = temp_mem[3297];
   memory[824][2] = temp_mem[3298];
   memory[824][3] = temp_mem[3299];

   memory[825][0] = temp_mem[3300];
   memory[825][1] = temp_mem[3301];
   memory[825][2] = temp_mem[3302];
   memory[825][3] = temp_mem[3303];

   memory[826][0] = temp_mem[3304];
   memory[826][1] = temp_mem[3305];
   memory[826][2] = temp_mem[3306];
   memory[826][3] = temp_mem[3307];

   memory[827][0] = temp_mem[3308];
   memory[827][1] = temp_mem[3309];
   memory[827][2] = temp_mem[3310];
   memory[827][3] = temp_mem[3311];

   memory[828][0] = temp_mem[3312];
   memory[828][1] = temp_mem[3313];
   memory[828][2] = temp_mem[3314];
   memory[828][3] = temp_mem[3315];

   memory[829][0] = temp_mem[3316];
   memory[829][1] = temp_mem[3317];
   memory[829][2] = temp_mem[3318];
   memory[829][3] = temp_mem[3319];

   memory[830][0] = temp_mem[3320];
   memory[830][1] = temp_mem[3321];
   memory[830][2] = temp_mem[3322];
   memory[830][3] = temp_mem[3323];

   memory[831][0] = temp_mem[3324];
   memory[831][1] = temp_mem[3325];
   memory[831][2] = temp_mem[3326];
   memory[831][3] = temp_mem[3327];

   memory[832][0] = temp_mem[3328];
   memory[832][1] = temp_mem[3329];
   memory[832][2] = temp_mem[3330];
   memory[832][3] = temp_mem[3331];

   memory[833][0] = temp_mem[3332];
   memory[833][1] = temp_mem[3333];
   memory[833][2] = temp_mem[3334];
   memory[833][3] = temp_mem[3335];

   memory[834][0] = temp_mem[3336];
   memory[834][1] = temp_mem[3337];
   memory[834][2] = temp_mem[3338];
   memory[834][3] = temp_mem[3339];

   memory[835][0] = temp_mem[3340];
   memory[835][1] = temp_mem[3341];
   memory[835][2] = temp_mem[3342];
   memory[835][3] = temp_mem[3343];

   memory[836][0] = temp_mem[3344];
   memory[836][1] = temp_mem[3345];
   memory[836][2] = temp_mem[3346];
   memory[836][3] = temp_mem[3347];

   memory[837][0] = temp_mem[3348];
   memory[837][1] = temp_mem[3349];
   memory[837][2] = temp_mem[3350];
   memory[837][3] = temp_mem[3351];

   memory[838][0] = temp_mem[3352];
   memory[838][1] = temp_mem[3353];
   memory[838][2] = temp_mem[3354];
   memory[838][3] = temp_mem[3355];

   memory[839][0] = temp_mem[3356];
   memory[839][1] = temp_mem[3357];
   memory[839][2] = temp_mem[3358];
   memory[839][3] = temp_mem[3359];

   memory[840][0] = temp_mem[3360];
   memory[840][1] = temp_mem[3361];
   memory[840][2] = temp_mem[3362];
   memory[840][3] = temp_mem[3363];

   memory[841][0] = temp_mem[3364];
   memory[841][1] = temp_mem[3365];
   memory[841][2] = temp_mem[3366];
   memory[841][3] = temp_mem[3367];

   memory[842][0] = temp_mem[3368];
   memory[842][1] = temp_mem[3369];
   memory[842][2] = temp_mem[3370];
   memory[842][3] = temp_mem[3371];

   memory[843][0] = temp_mem[3372];
   memory[843][1] = temp_mem[3373];
   memory[843][2] = temp_mem[3374];
   memory[843][3] = temp_mem[3375];

   memory[844][0] = temp_mem[3376];
   memory[844][1] = temp_mem[3377];
   memory[844][2] = temp_mem[3378];
   memory[844][3] = temp_mem[3379];

   memory[845][0] = temp_mem[3380];
   memory[845][1] = temp_mem[3381];
   memory[845][2] = temp_mem[3382];
   memory[845][3] = temp_mem[3383];

   memory[846][0] = temp_mem[3384];
   memory[846][1] = temp_mem[3385];
   memory[846][2] = temp_mem[3386];
   memory[846][3] = temp_mem[3387];

   memory[847][0] = temp_mem[3388];
   memory[847][1] = temp_mem[3389];
   memory[847][2] = temp_mem[3390];
   memory[847][3] = temp_mem[3391];

   memory[848][0] = temp_mem[3392];
   memory[848][1] = temp_mem[3393];
   memory[848][2] = temp_mem[3394];
   memory[848][3] = temp_mem[3395];

   memory[849][0] = temp_mem[3396];
   memory[849][1] = temp_mem[3397];
   memory[849][2] = temp_mem[3398];
   memory[849][3] = temp_mem[3399];

   memory[850][0] = temp_mem[3400];
   memory[850][1] = temp_mem[3401];
   memory[850][2] = temp_mem[3402];
   memory[850][3] = temp_mem[3403];

   memory[851][0] = temp_mem[3404];
   memory[851][1] = temp_mem[3405];
   memory[851][2] = temp_mem[3406];
   memory[851][3] = temp_mem[3407];

   memory[852][0] = temp_mem[3408];
   memory[852][1] = temp_mem[3409];
   memory[852][2] = temp_mem[3410];
   memory[852][3] = temp_mem[3411];

   memory[853][0] = temp_mem[3412];
   memory[853][1] = temp_mem[3413];
   memory[853][2] = temp_mem[3414];
   memory[853][3] = temp_mem[3415];

   memory[854][0] = temp_mem[3416];
   memory[854][1] = temp_mem[3417];
   memory[854][2] = temp_mem[3418];
   memory[854][3] = temp_mem[3419];

   memory[855][0] = temp_mem[3420];
   memory[855][1] = temp_mem[3421];
   memory[855][2] = temp_mem[3422];
   memory[855][3] = temp_mem[3423];

   memory[856][0] = temp_mem[3424];
   memory[856][1] = temp_mem[3425];
   memory[856][2] = temp_mem[3426];
   memory[856][3] = temp_mem[3427];

   memory[857][0] = temp_mem[3428];
   memory[857][1] = temp_mem[3429];
   memory[857][2] = temp_mem[3430];
   memory[857][3] = temp_mem[3431];

   memory[858][0] = temp_mem[3432];
   memory[858][1] = temp_mem[3433];
   memory[858][2] = temp_mem[3434];
   memory[858][3] = temp_mem[3435];

   memory[859][0] = temp_mem[3436];
   memory[859][1] = temp_mem[3437];
   memory[859][2] = temp_mem[3438];
   memory[859][3] = temp_mem[3439];

   memory[860][0] = temp_mem[3440];
   memory[860][1] = temp_mem[3441];
   memory[860][2] = temp_mem[3442];
   memory[860][3] = temp_mem[3443];

   memory[861][0] = temp_mem[3444];
   memory[861][1] = temp_mem[3445];
   memory[861][2] = temp_mem[3446];
   memory[861][3] = temp_mem[3447];

   memory[862][0] = temp_mem[3448];
   memory[862][1] = temp_mem[3449];
   memory[862][2] = temp_mem[3450];
   memory[862][3] = temp_mem[3451];

   memory[863][0] = temp_mem[3452];
   memory[863][1] = temp_mem[3453];
   memory[863][2] = temp_mem[3454];
   memory[863][3] = temp_mem[3455];

   memory[864][0] = temp_mem[3456];
   memory[864][1] = temp_mem[3457];
   memory[864][2] = temp_mem[3458];
   memory[864][3] = temp_mem[3459];

   memory[865][0] = temp_mem[3460];
   memory[865][1] = temp_mem[3461];
   memory[865][2] = temp_mem[3462];
   memory[865][3] = temp_mem[3463];

   memory[866][0] = temp_mem[3464];
   memory[866][1] = temp_mem[3465];
   memory[866][2] = temp_mem[3466];
   memory[866][3] = temp_mem[3467];

   memory[867][0] = temp_mem[3468];
   memory[867][1] = temp_mem[3469];
   memory[867][2] = temp_mem[3470];
   memory[867][3] = temp_mem[3471];

   memory[868][0] = temp_mem[3472];
   memory[868][1] = temp_mem[3473];
   memory[868][2] = temp_mem[3474];
   memory[868][3] = temp_mem[3475];

   memory[869][0] = temp_mem[3476];
   memory[869][1] = temp_mem[3477];
   memory[869][2] = temp_mem[3478];
   memory[869][3] = temp_mem[3479];

   memory[870][0] = temp_mem[3480];
   memory[870][1] = temp_mem[3481];
   memory[870][2] = temp_mem[3482];
   memory[870][3] = temp_mem[3483];

   memory[871][0] = temp_mem[3484];
   memory[871][1] = temp_mem[3485];
   memory[871][2] = temp_mem[3486];
   memory[871][3] = temp_mem[3487];

   memory[872][0] = temp_mem[3488];
   memory[872][1] = temp_mem[3489];
   memory[872][2] = temp_mem[3490];
   memory[872][3] = temp_mem[3491];

   memory[873][0] = temp_mem[3492];
   memory[873][1] = temp_mem[3493];
   memory[873][2] = temp_mem[3494];
   memory[873][3] = temp_mem[3495];

   memory[874][0] = temp_mem[3496];
   memory[874][1] = temp_mem[3497];
   memory[874][2] = temp_mem[3498];
   memory[874][3] = temp_mem[3499];

   memory[875][0] = temp_mem[3500];
   memory[875][1] = temp_mem[3501];
   memory[875][2] = temp_mem[3502];
   memory[875][3] = temp_mem[3503];

   memory[876][0] = temp_mem[3504];
   memory[876][1] = temp_mem[3505];
   memory[876][2] = temp_mem[3506];
   memory[876][3] = temp_mem[3507];

   memory[877][0] = temp_mem[3508];
   memory[877][1] = temp_mem[3509];
   memory[877][2] = temp_mem[3510];
   memory[877][3] = temp_mem[3511];

   memory[878][0] = temp_mem[3512];
   memory[878][1] = temp_mem[3513];
   memory[878][2] = temp_mem[3514];
   memory[878][3] = temp_mem[3515];

   memory[879][0] = temp_mem[3516];
   memory[879][1] = temp_mem[3517];
   memory[879][2] = temp_mem[3518];
   memory[879][3] = temp_mem[3519];

   memory[880][0] = temp_mem[3520];
   memory[880][1] = temp_mem[3521];
   memory[880][2] = temp_mem[3522];
   memory[880][3] = temp_mem[3523];

   memory[881][0] = temp_mem[3524];
   memory[881][1] = temp_mem[3525];
   memory[881][2] = temp_mem[3526];
   memory[881][3] = temp_mem[3527];

   memory[882][0] = temp_mem[3528];
   memory[882][1] = temp_mem[3529];
   memory[882][2] = temp_mem[3530];
   memory[882][3] = temp_mem[3531];

   memory[883][0] = temp_mem[3532];
   memory[883][1] = temp_mem[3533];
   memory[883][2] = temp_mem[3534];
   memory[883][3] = temp_mem[3535];

   memory[884][0] = temp_mem[3536];
   memory[884][1] = temp_mem[3537];
   memory[884][2] = temp_mem[3538];
   memory[884][3] = temp_mem[3539];

   memory[885][0] = temp_mem[3540];
   memory[885][1] = temp_mem[3541];
   memory[885][2] = temp_mem[3542];
   memory[885][3] = temp_mem[3543];

   memory[886][0] = temp_mem[3544];
   memory[886][1] = temp_mem[3545];
   memory[886][2] = temp_mem[3546];
   memory[886][3] = temp_mem[3547];

   memory[887][0] = temp_mem[3548];
   memory[887][1] = temp_mem[3549];
   memory[887][2] = temp_mem[3550];
   memory[887][3] = temp_mem[3551];

   memory[888][0] = temp_mem[3552];
   memory[888][1] = temp_mem[3553];
   memory[888][2] = temp_mem[3554];
   memory[888][3] = temp_mem[3555];

   memory[889][0] = temp_mem[3556];
   memory[889][1] = temp_mem[3557];
   memory[889][2] = temp_mem[3558];
   memory[889][3] = temp_mem[3559];

   memory[890][0] = temp_mem[3560];
   memory[890][1] = temp_mem[3561];
   memory[890][2] = temp_mem[3562];
   memory[890][3] = temp_mem[3563];

   memory[891][0] = temp_mem[3564];
   memory[891][1] = temp_mem[3565];
   memory[891][2] = temp_mem[3566];
   memory[891][3] = temp_mem[3567];

   memory[892][0] = temp_mem[3568];
   memory[892][1] = temp_mem[3569];
   memory[892][2] = temp_mem[3570];
   memory[892][3] = temp_mem[3571];

   memory[893][0] = temp_mem[3572];
   memory[893][1] = temp_mem[3573];
   memory[893][2] = temp_mem[3574];
   memory[893][3] = temp_mem[3575];

   memory[894][0] = temp_mem[3576];
   memory[894][1] = temp_mem[3577];
   memory[894][2] = temp_mem[3578];
   memory[894][3] = temp_mem[3579];

   memory[895][0] = temp_mem[3580];
   memory[895][1] = temp_mem[3581];
   memory[895][2] = temp_mem[3582];
   memory[895][3] = temp_mem[3583];

   memory[896][0] = temp_mem[3584];
   memory[896][1] = temp_mem[3585];
   memory[896][2] = temp_mem[3586];
   memory[896][3] = temp_mem[3587];

   memory[897][0] = temp_mem[3588];
   memory[897][1] = temp_mem[3589];
   memory[897][2] = temp_mem[3590];
   memory[897][3] = temp_mem[3591];

   memory[898][0] = temp_mem[3592];
   memory[898][1] = temp_mem[3593];
   memory[898][2] = temp_mem[3594];
   memory[898][3] = temp_mem[3595];

   memory[899][0] = temp_mem[3596];
   memory[899][1] = temp_mem[3597];
   memory[899][2] = temp_mem[3598];
   memory[899][3] = temp_mem[3599];

   memory[900][0] = temp_mem[3600];
   memory[900][1] = temp_mem[3601];
   memory[900][2] = temp_mem[3602];
   memory[900][3] = temp_mem[3603];

   memory[901][0] = temp_mem[3604];
   memory[901][1] = temp_mem[3605];
   memory[901][2] = temp_mem[3606];
   memory[901][3] = temp_mem[3607];

   memory[902][0] = temp_mem[3608];
   memory[902][1] = temp_mem[3609];
   memory[902][2] = temp_mem[3610];
   memory[902][3] = temp_mem[3611];

   memory[903][0] = temp_mem[3612];
   memory[903][1] = temp_mem[3613];
   memory[903][2] = temp_mem[3614];
   memory[903][3] = temp_mem[3615];

   memory[904][0] = temp_mem[3616];
   memory[904][1] = temp_mem[3617];
   memory[904][2] = temp_mem[3618];
   memory[904][3] = temp_mem[3619];

   memory[905][0] = temp_mem[3620];
   memory[905][1] = temp_mem[3621];
   memory[905][2] = temp_mem[3622];
   memory[905][3] = temp_mem[3623];

   memory[906][0] = temp_mem[3624];
   memory[906][1] = temp_mem[3625];
   memory[906][2] = temp_mem[3626];
   memory[906][3] = temp_mem[3627];

   memory[907][0] = temp_mem[3628];
   memory[907][1] = temp_mem[3629];
   memory[907][2] = temp_mem[3630];
   memory[907][3] = temp_mem[3631];

   memory[908][0] = temp_mem[3632];
   memory[908][1] = temp_mem[3633];
   memory[908][2] = temp_mem[3634];
   memory[908][3] = temp_mem[3635];

   memory[909][0] = temp_mem[3636];
   memory[909][1] = temp_mem[3637];
   memory[909][2] = temp_mem[3638];
   memory[909][3] = temp_mem[3639];

   memory[910][0] = temp_mem[3640];
   memory[910][1] = temp_mem[3641];
   memory[910][2] = temp_mem[3642];
   memory[910][3] = temp_mem[3643];

   memory[911][0] = temp_mem[3644];
   memory[911][1] = temp_mem[3645];
   memory[911][2] = temp_mem[3646];
   memory[911][3] = temp_mem[3647];

   memory[912][0] = temp_mem[3648];
   memory[912][1] = temp_mem[3649];
   memory[912][2] = temp_mem[3650];
   memory[912][3] = temp_mem[3651];

   memory[913][0] = temp_mem[3652];
   memory[913][1] = temp_mem[3653];
   memory[913][2] = temp_mem[3654];
   memory[913][3] = temp_mem[3655];

   memory[914][0] = temp_mem[3656];
   memory[914][1] = temp_mem[3657];
   memory[914][2] = temp_mem[3658];
   memory[914][3] = temp_mem[3659];

   memory[915][0] = temp_mem[3660];
   memory[915][1] = temp_mem[3661];
   memory[915][2] = temp_mem[3662];
   memory[915][3] = temp_mem[3663];

   memory[916][0] = temp_mem[3664];
   memory[916][1] = temp_mem[3665];
   memory[916][2] = temp_mem[3666];
   memory[916][3] = temp_mem[3667];

   memory[917][0] = temp_mem[3668];
   memory[917][1] = temp_mem[3669];
   memory[917][2] = temp_mem[3670];
   memory[917][3] = temp_mem[3671];

   memory[918][0] = temp_mem[3672];
   memory[918][1] = temp_mem[3673];
   memory[918][2] = temp_mem[3674];
   memory[918][3] = temp_mem[3675];

   memory[919][0] = temp_mem[3676];
   memory[919][1] = temp_mem[3677];
   memory[919][2] = temp_mem[3678];
   memory[919][3] = temp_mem[3679];

   memory[920][0] = temp_mem[3680];
   memory[920][1] = temp_mem[3681];
   memory[920][2] = temp_mem[3682];
   memory[920][3] = temp_mem[3683];

   memory[921][0] = temp_mem[3684];
   memory[921][1] = temp_mem[3685];
   memory[921][2] = temp_mem[3686];
   memory[921][3] = temp_mem[3687];

   memory[922][0] = temp_mem[3688];
   memory[922][1] = temp_mem[3689];
   memory[922][2] = temp_mem[3690];
   memory[922][3] = temp_mem[3691];

   memory[923][0] = temp_mem[3692];
   memory[923][1] = temp_mem[3693];
   memory[923][2] = temp_mem[3694];
   memory[923][3] = temp_mem[3695];

   memory[924][0] = temp_mem[3696];
   memory[924][1] = temp_mem[3697];
   memory[924][2] = temp_mem[3698];
   memory[924][3] = temp_mem[3699];

   memory[925][0] = temp_mem[3700];
   memory[925][1] = temp_mem[3701];
   memory[925][2] = temp_mem[3702];
   memory[925][3] = temp_mem[3703];

   memory[926][0] = temp_mem[3704];
   memory[926][1] = temp_mem[3705];
   memory[926][2] = temp_mem[3706];
   memory[926][3] = temp_mem[3707];

   memory[927][0] = temp_mem[3708];
   memory[927][1] = temp_mem[3709];
   memory[927][2] = temp_mem[3710];
   memory[927][3] = temp_mem[3711];

   memory[928][0] = temp_mem[3712];
   memory[928][1] = temp_mem[3713];
   memory[928][2] = temp_mem[3714];
   memory[928][3] = temp_mem[3715];

   memory[929][0] = temp_mem[3716];
   memory[929][1] = temp_mem[3717];
   memory[929][2] = temp_mem[3718];
   memory[929][3] = temp_mem[3719];

   memory[930][0] = temp_mem[3720];
   memory[930][1] = temp_mem[3721];
   memory[930][2] = temp_mem[3722];
   memory[930][3] = temp_mem[3723];

   memory[931][0] = temp_mem[3724];
   memory[931][1] = temp_mem[3725];
   memory[931][2] = temp_mem[3726];
   memory[931][3] = temp_mem[3727];

   memory[932][0] = temp_mem[3728];
   memory[932][1] = temp_mem[3729];
   memory[932][2] = temp_mem[3730];
   memory[932][3] = temp_mem[3731];

   memory[933][0] = temp_mem[3732];
   memory[933][1] = temp_mem[3733];
   memory[933][2] = temp_mem[3734];
   memory[933][3] = temp_mem[3735];

   memory[934][0] = temp_mem[3736];
   memory[934][1] = temp_mem[3737];
   memory[934][2] = temp_mem[3738];
   memory[934][3] = temp_mem[3739];

   memory[935][0] = temp_mem[3740];
   memory[935][1] = temp_mem[3741];
   memory[935][2] = temp_mem[3742];
   memory[935][3] = temp_mem[3743];

   memory[936][0] = temp_mem[3744];
   memory[936][1] = temp_mem[3745];
   memory[936][2] = temp_mem[3746];
   memory[936][3] = temp_mem[3747];

   memory[937][0] = temp_mem[3748];
   memory[937][1] = temp_mem[3749];
   memory[937][2] = temp_mem[3750];
   memory[937][3] = temp_mem[3751];

   memory[938][0] = temp_mem[3752];
   memory[938][1] = temp_mem[3753];
   memory[938][2] = temp_mem[3754];
   memory[938][3] = temp_mem[3755];

   memory[939][0] = temp_mem[3756];
   memory[939][1] = temp_mem[3757];
   memory[939][2] = temp_mem[3758];
   memory[939][3] = temp_mem[3759];

   memory[940][0] = temp_mem[3760];
   memory[940][1] = temp_mem[3761];
   memory[940][2] = temp_mem[3762];
   memory[940][3] = temp_mem[3763];

   memory[941][0] = temp_mem[3764];
   memory[941][1] = temp_mem[3765];
   memory[941][2] = temp_mem[3766];
   memory[941][3] = temp_mem[3767];

   memory[942][0] = temp_mem[3768];
   memory[942][1] = temp_mem[3769];
   memory[942][2] = temp_mem[3770];
   memory[942][3] = temp_mem[3771];

   memory[943][0] = temp_mem[3772];
   memory[943][1] = temp_mem[3773];
   memory[943][2] = temp_mem[3774];
   memory[943][3] = temp_mem[3775];

   memory[944][0] = temp_mem[3776];
   memory[944][1] = temp_mem[3777];
   memory[944][2] = temp_mem[3778];
   memory[944][3] = temp_mem[3779];

   memory[945][0] = temp_mem[3780];
   memory[945][1] = temp_mem[3781];
   memory[945][2] = temp_mem[3782];
   memory[945][3] = temp_mem[3783];

   memory[946][0] = temp_mem[3784];
   memory[946][1] = temp_mem[3785];
   memory[946][2] = temp_mem[3786];
   memory[946][3] = temp_mem[3787];

   memory[947][0] = temp_mem[3788];
   memory[947][1] = temp_mem[3789];
   memory[947][2] = temp_mem[3790];
   memory[947][3] = temp_mem[3791];

   memory[948][0] = temp_mem[3792];
   memory[948][1] = temp_mem[3793];
   memory[948][2] = temp_mem[3794];
   memory[948][3] = temp_mem[3795];

   memory[949][0] = temp_mem[3796];
   memory[949][1] = temp_mem[3797];
   memory[949][2] = temp_mem[3798];
   memory[949][3] = temp_mem[3799];

   memory[950][0] = temp_mem[3800];
   memory[950][1] = temp_mem[3801];
   memory[950][2] = temp_mem[3802];
   memory[950][3] = temp_mem[3803];

   memory[951][0] = temp_mem[3804];
   memory[951][1] = temp_mem[3805];
   memory[951][2] = temp_mem[3806];
   memory[951][3] = temp_mem[3807];

   memory[952][0] = temp_mem[3808];
   memory[952][1] = temp_mem[3809];
   memory[952][2] = temp_mem[3810];
   memory[952][3] = temp_mem[3811];

   memory[953][0] = temp_mem[3812];
   memory[953][1] = temp_mem[3813];
   memory[953][2] = temp_mem[3814];
   memory[953][3] = temp_mem[3815];

   memory[954][0] = temp_mem[3816];
   memory[954][1] = temp_mem[3817];
   memory[954][2] = temp_mem[3818];
   memory[954][3] = temp_mem[3819];

   memory[955][0] = temp_mem[3820];
   memory[955][1] = temp_mem[3821];
   memory[955][2] = temp_mem[3822];
   memory[955][3] = temp_mem[3823];

   memory[956][0] = temp_mem[3824];
   memory[956][1] = temp_mem[3825];
   memory[956][2] = temp_mem[3826];
   memory[956][3] = temp_mem[3827];

   memory[957][0] = temp_mem[3828];
   memory[957][1] = temp_mem[3829];
   memory[957][2] = temp_mem[3830];
   memory[957][3] = temp_mem[3831];

   memory[958][0] = temp_mem[3832];
   memory[958][1] = temp_mem[3833];
   memory[958][2] = temp_mem[3834];
   memory[958][3] = temp_mem[3835];

   memory[959][0] = temp_mem[3836];
   memory[959][1] = temp_mem[3837];
   memory[959][2] = temp_mem[3838];
   memory[959][3] = temp_mem[3839];

   memory[960][0] = temp_mem[3840];
   memory[960][1] = temp_mem[3841];
   memory[960][2] = temp_mem[3842];
   memory[960][3] = temp_mem[3843];

   memory[961][0] = temp_mem[3844];
   memory[961][1] = temp_mem[3845];
   memory[961][2] = temp_mem[3846];
   memory[961][3] = temp_mem[3847];

   memory[962][0] = temp_mem[3848];
   memory[962][1] = temp_mem[3849];
   memory[962][2] = temp_mem[3850];
   memory[962][3] = temp_mem[3851];

   memory[963][0] = temp_mem[3852];
   memory[963][1] = temp_mem[3853];
   memory[963][2] = temp_mem[3854];
   memory[963][3] = temp_mem[3855];

   memory[964][0] = temp_mem[3856];
   memory[964][1] = temp_mem[3857];
   memory[964][2] = temp_mem[3858];
   memory[964][3] = temp_mem[3859];

   memory[965][0] = temp_mem[3860];
   memory[965][1] = temp_mem[3861];
   memory[965][2] = temp_mem[3862];
   memory[965][3] = temp_mem[3863];

   memory[966][0] = temp_mem[3864];
   memory[966][1] = temp_mem[3865];
   memory[966][2] = temp_mem[3866];
   memory[966][3] = temp_mem[3867];

   memory[967][0] = temp_mem[3868];
   memory[967][1] = temp_mem[3869];
   memory[967][2] = temp_mem[3870];
   memory[967][3] = temp_mem[3871];

   memory[968][0] = temp_mem[3872];
   memory[968][1] = temp_mem[3873];
   memory[968][2] = temp_mem[3874];
   memory[968][3] = temp_mem[3875];

   memory[969][0] = temp_mem[3876];
   memory[969][1] = temp_mem[3877];
   memory[969][2] = temp_mem[3878];
   memory[969][3] = temp_mem[3879];

   memory[970][0] = temp_mem[3880];
   memory[970][1] = temp_mem[3881];
   memory[970][2] = temp_mem[3882];
   memory[970][3] = temp_mem[3883];

   memory[971][0] = temp_mem[3884];
   memory[971][1] = temp_mem[3885];
   memory[971][2] = temp_mem[3886];
   memory[971][3] = temp_mem[3887];

   memory[972][0] = temp_mem[3888];
   memory[972][1] = temp_mem[3889];
   memory[972][2] = temp_mem[3890];
   memory[972][3] = temp_mem[3891];

   memory[973][0] = temp_mem[3892];
   memory[973][1] = temp_mem[3893];
   memory[973][2] = temp_mem[3894];
   memory[973][3] = temp_mem[3895];

   memory[974][0] = temp_mem[3896];
   memory[974][1] = temp_mem[3897];
   memory[974][2] = temp_mem[3898];
   memory[974][3] = temp_mem[3899];

   memory[975][0] = temp_mem[3900];
   memory[975][1] = temp_mem[3901];
   memory[975][2] = temp_mem[3902];
   memory[975][3] = temp_mem[3903];

   memory[976][0] = temp_mem[3904];
   memory[976][1] = temp_mem[3905];
   memory[976][2] = temp_mem[3906];
   memory[976][3] = temp_mem[3907];

   memory[977][0] = temp_mem[3908];
   memory[977][1] = temp_mem[3909];
   memory[977][2] = temp_mem[3910];
   memory[977][3] = temp_mem[3911];

   memory[978][0] = temp_mem[3912];
   memory[978][1] = temp_mem[3913];
   memory[978][2] = temp_mem[3914];
   memory[978][3] = temp_mem[3915];

   memory[979][0] = temp_mem[3916];
   memory[979][1] = temp_mem[3917];
   memory[979][2] = temp_mem[3918];
   memory[979][3] = temp_mem[3919];

   memory[980][0] = temp_mem[3920];
   memory[980][1] = temp_mem[3921];
   memory[980][2] = temp_mem[3922];
   memory[980][3] = temp_mem[3923];

   memory[981][0] = temp_mem[3924];
   memory[981][1] = temp_mem[3925];
   memory[981][2] = temp_mem[3926];
   memory[981][3] = temp_mem[3927];

   memory[982][0] = temp_mem[3928];
   memory[982][1] = temp_mem[3929];
   memory[982][2] = temp_mem[3930];
   memory[982][3] = temp_mem[3931];

   memory[983][0] = temp_mem[3932];
   memory[983][1] = temp_mem[3933];
   memory[983][2] = temp_mem[3934];
   memory[983][3] = temp_mem[3935];

   memory[984][0] = temp_mem[3936];
   memory[984][1] = temp_mem[3937];
   memory[984][2] = temp_mem[3938];
   memory[984][3] = temp_mem[3939];

   memory[985][0] = temp_mem[3940];
   memory[985][1] = temp_mem[3941];
   memory[985][2] = temp_mem[3942];
   memory[985][3] = temp_mem[3943];

   memory[986][0] = temp_mem[3944];
   memory[986][1] = temp_mem[3945];
   memory[986][2] = temp_mem[3946];
   memory[986][3] = temp_mem[3947];

   memory[987][0] = temp_mem[3948];
   memory[987][1] = temp_mem[3949];
   memory[987][2] = temp_mem[3950];
   memory[987][3] = temp_mem[3951];

   memory[988][0] = temp_mem[3952];
   memory[988][1] = temp_mem[3953];
   memory[988][2] = temp_mem[3954];
   memory[988][3] = temp_mem[3955];

   memory[989][0] = temp_mem[3956];
   memory[989][1] = temp_mem[3957];
   memory[989][2] = temp_mem[3958];
   memory[989][3] = temp_mem[3959];

   memory[990][0] = temp_mem[3960];
   memory[990][1] = temp_mem[3961];
   memory[990][2] = temp_mem[3962];
   memory[990][3] = temp_mem[3963];

   memory[991][0] = temp_mem[3964];
   memory[991][1] = temp_mem[3965];
   memory[991][2] = temp_mem[3966];
   memory[991][3] = temp_mem[3967];

   memory[992][0] = temp_mem[3968];
   memory[992][1] = temp_mem[3969];
   memory[992][2] = temp_mem[3970];
   memory[992][3] = temp_mem[3971];

   memory[993][0] = temp_mem[3972];
   memory[993][1] = temp_mem[3973];
   memory[993][2] = temp_mem[3974];
   memory[993][3] = temp_mem[3975];

   memory[994][0] = temp_mem[3976];
   memory[994][1] = temp_mem[3977];
   memory[994][2] = temp_mem[3978];
   memory[994][3] = temp_mem[3979];

   memory[995][0] = temp_mem[3980];
   memory[995][1] = temp_mem[3981];
   memory[995][2] = temp_mem[3982];
   memory[995][3] = temp_mem[3983];

   memory[996][0] = temp_mem[3984];
   memory[996][1] = temp_mem[3985];
   memory[996][2] = temp_mem[3986];
   memory[996][3] = temp_mem[3987];

   memory[997][0] = temp_mem[3988];
   memory[997][1] = temp_mem[3989];
   memory[997][2] = temp_mem[3990];
   memory[997][3] = temp_mem[3991];

   memory[998][0] = temp_mem[3992];
   memory[998][1] = temp_mem[3993];
   memory[998][2] = temp_mem[3994];
   memory[998][3] = temp_mem[3995];

   memory[999][0] = temp_mem[3996];
   memory[999][1] = temp_mem[3997];
   memory[999][2] = temp_mem[3998];
   memory[999][3] = temp_mem[3999];

   memory[1000][0] = temp_mem[4000];
   memory[1000][1] = temp_mem[4001];
   memory[1000][2] = temp_mem[4002];
   memory[1000][3] = temp_mem[4003];

   memory[1001][0] = temp_mem[4004];
   memory[1001][1] = temp_mem[4005];
   memory[1001][2] = temp_mem[4006];
   memory[1001][3] = temp_mem[4007];

   memory[1002][0] = temp_mem[4008];
   memory[1002][1] = temp_mem[4009];
   memory[1002][2] = temp_mem[4010];
   memory[1002][3] = temp_mem[4011];

   memory[1003][0] = temp_mem[4012];
   memory[1003][1] = temp_mem[4013];
   memory[1003][2] = temp_mem[4014];
   memory[1003][3] = temp_mem[4015];

   memory[1004][0] = temp_mem[4016];
   memory[1004][1] = temp_mem[4017];
   memory[1004][2] = temp_mem[4018];
   memory[1004][3] = temp_mem[4019];

   memory[1005][0] = temp_mem[4020];
   memory[1005][1] = temp_mem[4021];
   memory[1005][2] = temp_mem[4022];
   memory[1005][3] = temp_mem[4023];

   memory[1006][0] = temp_mem[4024];
   memory[1006][1] = temp_mem[4025];
   memory[1006][2] = temp_mem[4026];
   memory[1006][3] = temp_mem[4027];

   memory[1007][0] = temp_mem[4028];
   memory[1007][1] = temp_mem[4029];
   memory[1007][2] = temp_mem[4030];
   memory[1007][3] = temp_mem[4031];

   memory[1008][0] = temp_mem[4032];
   memory[1008][1] = temp_mem[4033];
   memory[1008][2] = temp_mem[4034];
   memory[1008][3] = temp_mem[4035];

   memory[1009][0] = temp_mem[4036];
   memory[1009][1] = temp_mem[4037];
   memory[1009][2] = temp_mem[4038];
   memory[1009][3] = temp_mem[4039];

   memory[1010][0] = temp_mem[4040];
   memory[1010][1] = temp_mem[4041];
   memory[1010][2] = temp_mem[4042];
   memory[1010][3] = temp_mem[4043];

   memory[1011][0] = temp_mem[4044];
   memory[1011][1] = temp_mem[4045];
   memory[1011][2] = temp_mem[4046];
   memory[1011][3] = temp_mem[4047];

   memory[1012][0] = temp_mem[4048];
   memory[1012][1] = temp_mem[4049];
   memory[1012][2] = temp_mem[4050];
   memory[1012][3] = temp_mem[4051];

   memory[1013][0] = temp_mem[4052];
   memory[1013][1] = temp_mem[4053];
   memory[1013][2] = temp_mem[4054];
   memory[1013][3] = temp_mem[4055];

   memory[1014][0] = temp_mem[4056];
   memory[1014][1] = temp_mem[4057];
   memory[1014][2] = temp_mem[4058];
   memory[1014][3] = temp_mem[4059];

   memory[1015][0] = temp_mem[4060];
   memory[1015][1] = temp_mem[4061];
   memory[1015][2] = temp_mem[4062];
   memory[1015][3] = temp_mem[4063];

   memory[1016][0] = temp_mem[4064];
   memory[1016][1] = temp_mem[4065];
   memory[1016][2] = temp_mem[4066];
   memory[1016][3] = temp_mem[4067];

   memory[1017][0] = temp_mem[4068];
   memory[1017][1] = temp_mem[4069];
   memory[1017][2] = temp_mem[4070];
   memory[1017][3] = temp_mem[4071];

   memory[1018][0] = temp_mem[4072];
   memory[1018][1] = temp_mem[4073];
   memory[1018][2] = temp_mem[4074];
   memory[1018][3] = temp_mem[4075];

   memory[1019][0] = temp_mem[4076];
   memory[1019][1] = temp_mem[4077];
   memory[1019][2] = temp_mem[4078];
   memory[1019][3] = temp_mem[4079];

   memory[1020][0] = temp_mem[4080];
   memory[1020][1] = temp_mem[4081];
   memory[1020][2] = temp_mem[4082];
   memory[1020][3] = temp_mem[4083];

   memory[1021][0] = temp_mem[4084];
   memory[1021][1] = temp_mem[4085];
   memory[1021][2] = temp_mem[4086];
   memory[1021][3] = temp_mem[4087];

   memory[1022][0] = temp_mem[4088];
   memory[1022][1] = temp_mem[4089];
   memory[1022][2] = temp_mem[4090];
   memory[1022][3] = temp_mem[4091];

   memory[1023][0] = temp_mem[4092];
   memory[1023][1] = temp_mem[4093];
   memory[1023][2] = temp_mem[4094];
   memory[1023][3] = temp_mem[4095];

   memory[1024][0] = temp_mem[4096];
   memory[1024][1] = temp_mem[4097];
   memory[1024][2] = temp_mem[4098];
   memory[1024][3] = temp_mem[4099];

   memory[1025][0] = temp_mem[4100];
   memory[1025][1] = temp_mem[4101];
   memory[1025][2] = temp_mem[4102];
   memory[1025][3] = temp_mem[4103];

   memory[1026][0] = temp_mem[4104];
   memory[1026][1] = temp_mem[4105];
   memory[1026][2] = temp_mem[4106];
   memory[1026][3] = temp_mem[4107];

   memory[1027][0] = temp_mem[4108];
   memory[1027][1] = temp_mem[4109];
   memory[1027][2] = temp_mem[4110];
   memory[1027][3] = temp_mem[4111];

   memory[1028][0] = temp_mem[4112];
   memory[1028][1] = temp_mem[4113];
   memory[1028][2] = temp_mem[4114];
   memory[1028][3] = temp_mem[4115];

   memory[1029][0] = temp_mem[4116];
   memory[1029][1] = temp_mem[4117];
   memory[1029][2] = temp_mem[4118];
   memory[1029][3] = temp_mem[4119];

   memory[1030][0] = temp_mem[4120];
   memory[1030][1] = temp_mem[4121];
   memory[1030][2] = temp_mem[4122];
   memory[1030][3] = temp_mem[4123];

   memory[1031][0] = temp_mem[4124];
   memory[1031][1] = temp_mem[4125];
   memory[1031][2] = temp_mem[4126];
   memory[1031][3] = temp_mem[4127];

   memory[1032][0] = temp_mem[4128];
   memory[1032][1] = temp_mem[4129];
   memory[1032][2] = temp_mem[4130];
   memory[1032][3] = temp_mem[4131];

   memory[1033][0] = temp_mem[4132];
   memory[1033][1] = temp_mem[4133];
   memory[1033][2] = temp_mem[4134];
   memory[1033][3] = temp_mem[4135];

   memory[1034][0] = temp_mem[4136];
   memory[1034][1] = temp_mem[4137];
   memory[1034][2] = temp_mem[4138];
   memory[1034][3] = temp_mem[4139];

   memory[1035][0] = temp_mem[4140];
   memory[1035][1] = temp_mem[4141];
   memory[1035][2] = temp_mem[4142];
   memory[1035][3] = temp_mem[4143];

   memory[1036][0] = temp_mem[4144];
   memory[1036][1] = temp_mem[4145];
   memory[1036][2] = temp_mem[4146];
   memory[1036][3] = temp_mem[4147];

   memory[1037][0] = temp_mem[4148];
   memory[1037][1] = temp_mem[4149];
   memory[1037][2] = temp_mem[4150];
   memory[1037][3] = temp_mem[4151];

   memory[1038][0] = temp_mem[4152];
   memory[1038][1] = temp_mem[4153];
   memory[1038][2] = temp_mem[4154];
   memory[1038][3] = temp_mem[4155];

   memory[1039][0] = temp_mem[4156];
   memory[1039][1] = temp_mem[4157];
   memory[1039][2] = temp_mem[4158];
   memory[1039][3] = temp_mem[4159];

   memory[1040][0] = temp_mem[4160];
   memory[1040][1] = temp_mem[4161];
   memory[1040][2] = temp_mem[4162];
   memory[1040][3] = temp_mem[4163];

   memory[1041][0] = temp_mem[4164];
   memory[1041][1] = temp_mem[4165];
   memory[1041][2] = temp_mem[4166];
   memory[1041][3] = temp_mem[4167];

   memory[1042][0] = temp_mem[4168];
   memory[1042][1] = temp_mem[4169];
   memory[1042][2] = temp_mem[4170];
   memory[1042][3] = temp_mem[4171];

   memory[1043][0] = temp_mem[4172];
   memory[1043][1] = temp_mem[4173];
   memory[1043][2] = temp_mem[4174];
   memory[1043][3] = temp_mem[4175];

   memory[1044][0] = temp_mem[4176];
   memory[1044][1] = temp_mem[4177];
   memory[1044][2] = temp_mem[4178];
   memory[1044][3] = temp_mem[4179];

   memory[1045][0] = temp_mem[4180];
   memory[1045][1] = temp_mem[4181];
   memory[1045][2] = temp_mem[4182];
   memory[1045][3] = temp_mem[4183];

   memory[1046][0] = temp_mem[4184];
   memory[1046][1] = temp_mem[4185];
   memory[1046][2] = temp_mem[4186];
   memory[1046][3] = temp_mem[4187];

   memory[1047][0] = temp_mem[4188];
   memory[1047][1] = temp_mem[4189];
   memory[1047][2] = temp_mem[4190];
   memory[1047][3] = temp_mem[4191];

   memory[1048][0] = temp_mem[4192];
   memory[1048][1] = temp_mem[4193];
   memory[1048][2] = temp_mem[4194];
   memory[1048][3] = temp_mem[4195];

   memory[1049][0] = temp_mem[4196];
   memory[1049][1] = temp_mem[4197];
   memory[1049][2] = temp_mem[4198];
   memory[1049][3] = temp_mem[4199];

   memory[1050][0] = temp_mem[4200];
   memory[1050][1] = temp_mem[4201];
   memory[1050][2] = temp_mem[4202];
   memory[1050][3] = temp_mem[4203];

   memory[1051][0] = temp_mem[4204];
   memory[1051][1] = temp_mem[4205];
   memory[1051][2] = temp_mem[4206];
   memory[1051][3] = temp_mem[4207];

   memory[1052][0] = temp_mem[4208];
   memory[1052][1] = temp_mem[4209];
   memory[1052][2] = temp_mem[4210];
   memory[1052][3] = temp_mem[4211];

   memory[1053][0] = temp_mem[4212];
   memory[1053][1] = temp_mem[4213];
   memory[1053][2] = temp_mem[4214];
   memory[1053][3] = temp_mem[4215];

   memory[1054][0] = temp_mem[4216];
   memory[1054][1] = temp_mem[4217];
   memory[1054][2] = temp_mem[4218];
   memory[1054][3] = temp_mem[4219];

   memory[1055][0] = temp_mem[4220];
   memory[1055][1] = temp_mem[4221];
   memory[1055][2] = temp_mem[4222];
   memory[1055][3] = temp_mem[4223];

   memory[1056][0] = temp_mem[4224];
   memory[1056][1] = temp_mem[4225];
   memory[1056][2] = temp_mem[4226];
   memory[1056][3] = temp_mem[4227];

   memory[1057][0] = temp_mem[4228];
   memory[1057][1] = temp_mem[4229];
   memory[1057][2] = temp_mem[4230];
   memory[1057][3] = temp_mem[4231];

   memory[1058][0] = temp_mem[4232];
   memory[1058][1] = temp_mem[4233];
   memory[1058][2] = temp_mem[4234];
   memory[1058][3] = temp_mem[4235];

   memory[1059][0] = temp_mem[4236];
   memory[1059][1] = temp_mem[4237];
   memory[1059][2] = temp_mem[4238];
   memory[1059][3] = temp_mem[4239];

   memory[1060][0] = temp_mem[4240];
   memory[1060][1] = temp_mem[4241];
   memory[1060][2] = temp_mem[4242];
   memory[1060][3] = temp_mem[4243];

   memory[1061][0] = temp_mem[4244];
   memory[1061][1] = temp_mem[4245];
   memory[1061][2] = temp_mem[4246];
   memory[1061][3] = temp_mem[4247];

   memory[1062][0] = temp_mem[4248];
   memory[1062][1] = temp_mem[4249];
   memory[1062][2] = temp_mem[4250];
   memory[1062][3] = temp_mem[4251];

   memory[1063][0] = temp_mem[4252];
   memory[1063][1] = temp_mem[4253];
   memory[1063][2] = temp_mem[4254];
   memory[1063][3] = temp_mem[4255];

   memory[1064][0] = temp_mem[4256];
   memory[1064][1] = temp_mem[4257];
   memory[1064][2] = temp_mem[4258];
   memory[1064][3] = temp_mem[4259];

   memory[1065][0] = temp_mem[4260];
   memory[1065][1] = temp_mem[4261];
   memory[1065][2] = temp_mem[4262];
   memory[1065][3] = temp_mem[4263];

   memory[1066][0] = temp_mem[4264];
   memory[1066][1] = temp_mem[4265];
   memory[1066][2] = temp_mem[4266];
   memory[1066][3] = temp_mem[4267];

   memory[1067][0] = temp_mem[4268];
   memory[1067][1] = temp_mem[4269];
   memory[1067][2] = temp_mem[4270];
   memory[1067][3] = temp_mem[4271];

   memory[1068][0] = temp_mem[4272];
   memory[1068][1] = temp_mem[4273];
   memory[1068][2] = temp_mem[4274];
   memory[1068][3] = temp_mem[4275];

   memory[1069][0] = temp_mem[4276];
   memory[1069][1] = temp_mem[4277];
   memory[1069][2] = temp_mem[4278];
   memory[1069][3] = temp_mem[4279];

   memory[1070][0] = temp_mem[4280];
   memory[1070][1] = temp_mem[4281];
   memory[1070][2] = temp_mem[4282];
   memory[1070][3] = temp_mem[4283];

   memory[1071][0] = temp_mem[4284];
   memory[1071][1] = temp_mem[4285];
   memory[1071][2] = temp_mem[4286];
   memory[1071][3] = temp_mem[4287];

   memory[1072][0] = temp_mem[4288];
   memory[1072][1] = temp_mem[4289];
   memory[1072][2] = temp_mem[4290];
   memory[1072][3] = temp_mem[4291];

   memory[1073][0] = temp_mem[4292];
   memory[1073][1] = temp_mem[4293];
   memory[1073][2] = temp_mem[4294];
   memory[1073][3] = temp_mem[4295];

   memory[1074][0] = temp_mem[4296];
   memory[1074][1] = temp_mem[4297];
   memory[1074][2] = temp_mem[4298];
   memory[1074][3] = temp_mem[4299];

   memory[1075][0] = temp_mem[4300];
   memory[1075][1] = temp_mem[4301];
   memory[1075][2] = temp_mem[4302];
   memory[1075][3] = temp_mem[4303];

   memory[1076][0] = temp_mem[4304];
   memory[1076][1] = temp_mem[4305];
   memory[1076][2] = temp_mem[4306];
   memory[1076][3] = temp_mem[4307];

   memory[1077][0] = temp_mem[4308];
   memory[1077][1] = temp_mem[4309];
   memory[1077][2] = temp_mem[4310];
   memory[1077][3] = temp_mem[4311];

   memory[1078][0] = temp_mem[4312];
   memory[1078][1] = temp_mem[4313];
   memory[1078][2] = temp_mem[4314];
   memory[1078][3] = temp_mem[4315];

   memory[1079][0] = temp_mem[4316];
   memory[1079][1] = temp_mem[4317];
   memory[1079][2] = temp_mem[4318];
   memory[1079][3] = temp_mem[4319];

   memory[1080][0] = temp_mem[4320];
   memory[1080][1] = temp_mem[4321];
   memory[1080][2] = temp_mem[4322];
   memory[1080][3] = temp_mem[4323];

   memory[1081][0] = temp_mem[4324];
   memory[1081][1] = temp_mem[4325];
   memory[1081][2] = temp_mem[4326];
   memory[1081][3] = temp_mem[4327];

   memory[1082][0] = temp_mem[4328];
   memory[1082][1] = temp_mem[4329];
   memory[1082][2] = temp_mem[4330];
   memory[1082][3] = temp_mem[4331];

   memory[1083][0] = temp_mem[4332];
   memory[1083][1] = temp_mem[4333];
   memory[1083][2] = temp_mem[4334];
   memory[1083][3] = temp_mem[4335];

   memory[1084][0] = temp_mem[4336];
   memory[1084][1] = temp_mem[4337];
   memory[1084][2] = temp_mem[4338];
   memory[1084][3] = temp_mem[4339];

   memory[1085][0] = temp_mem[4340];
   memory[1085][1] = temp_mem[4341];
   memory[1085][2] = temp_mem[4342];
   memory[1085][3] = temp_mem[4343];

   memory[1086][0] = temp_mem[4344];
   memory[1086][1] = temp_mem[4345];
   memory[1086][2] = temp_mem[4346];
   memory[1086][3] = temp_mem[4347];

   memory[1087][0] = temp_mem[4348];
   memory[1087][1] = temp_mem[4349];
   memory[1087][2] = temp_mem[4350];
   memory[1087][3] = temp_mem[4351];

   memory[1088][0] = temp_mem[4352];
   memory[1088][1] = temp_mem[4353];
   memory[1088][2] = temp_mem[4354];
   memory[1088][3] = temp_mem[4355];

   memory[1089][0] = temp_mem[4356];
   memory[1089][1] = temp_mem[4357];
   memory[1089][2] = temp_mem[4358];
   memory[1089][3] = temp_mem[4359];

   memory[1090][0] = temp_mem[4360];
   memory[1090][1] = temp_mem[4361];
   memory[1090][2] = temp_mem[4362];
   memory[1090][3] = temp_mem[4363];

   memory[1091][0] = temp_mem[4364];
   memory[1091][1] = temp_mem[4365];
   memory[1091][2] = temp_mem[4366];
   memory[1091][3] = temp_mem[4367];

   memory[1092][0] = temp_mem[4368];
   memory[1092][1] = temp_mem[4369];
   memory[1092][2] = temp_mem[4370];
   memory[1092][3] = temp_mem[4371];

   memory[1093][0] = temp_mem[4372];
   memory[1093][1] = temp_mem[4373];
   memory[1093][2] = temp_mem[4374];
   memory[1093][3] = temp_mem[4375];

   memory[1094][0] = temp_mem[4376];
   memory[1094][1] = temp_mem[4377];
   memory[1094][2] = temp_mem[4378];
   memory[1094][3] = temp_mem[4379];

   memory[1095][0] = temp_mem[4380];
   memory[1095][1] = temp_mem[4381];
   memory[1095][2] = temp_mem[4382];
   memory[1095][3] = temp_mem[4383];

   memory[1096][0] = temp_mem[4384];
   memory[1096][1] = temp_mem[4385];
   memory[1096][2] = temp_mem[4386];
   memory[1096][3] = temp_mem[4387];

   memory[1097][0] = temp_mem[4388];
   memory[1097][1] = temp_mem[4389];
   memory[1097][2] = temp_mem[4390];
   memory[1097][3] = temp_mem[4391];

   memory[1098][0] = temp_mem[4392];
   memory[1098][1] = temp_mem[4393];
   memory[1098][2] = temp_mem[4394];
   memory[1098][3] = temp_mem[4395];

   memory[1099][0] = temp_mem[4396];
   memory[1099][1] = temp_mem[4397];
   memory[1099][2] = temp_mem[4398];
   memory[1099][3] = temp_mem[4399];

   memory[1100][0] = temp_mem[4400];
   memory[1100][1] = temp_mem[4401];
   memory[1100][2] = temp_mem[4402];
   memory[1100][3] = temp_mem[4403];

   memory[1101][0] = temp_mem[4404];
   memory[1101][1] = temp_mem[4405];
   memory[1101][2] = temp_mem[4406];
   memory[1101][3] = temp_mem[4407];

   memory[1102][0] = temp_mem[4408];
   memory[1102][1] = temp_mem[4409];
   memory[1102][2] = temp_mem[4410];
   memory[1102][3] = temp_mem[4411];

   memory[1103][0] = temp_mem[4412];
   memory[1103][1] = temp_mem[4413];
   memory[1103][2] = temp_mem[4414];
   memory[1103][3] = temp_mem[4415];

   memory[1104][0] = temp_mem[4416];
   memory[1104][1] = temp_mem[4417];
   memory[1104][2] = temp_mem[4418];
   memory[1104][3] = temp_mem[4419];

   memory[1105][0] = temp_mem[4420];
   memory[1105][1] = temp_mem[4421];
   memory[1105][2] = temp_mem[4422];
   memory[1105][3] = temp_mem[4423];

   memory[1106][0] = temp_mem[4424];
   memory[1106][1] = temp_mem[4425];
   memory[1106][2] = temp_mem[4426];
   memory[1106][3] = temp_mem[4427];

   memory[1107][0] = temp_mem[4428];
   memory[1107][1] = temp_mem[4429];
   memory[1107][2] = temp_mem[4430];
   memory[1107][3] = temp_mem[4431];

   memory[1108][0] = temp_mem[4432];
   memory[1108][1] = temp_mem[4433];
   memory[1108][2] = temp_mem[4434];
   memory[1108][3] = temp_mem[4435];

   memory[1109][0] = temp_mem[4436];
   memory[1109][1] = temp_mem[4437];
   memory[1109][2] = temp_mem[4438];
   memory[1109][3] = temp_mem[4439];

   memory[1110][0] = temp_mem[4440];
   memory[1110][1] = temp_mem[4441];
   memory[1110][2] = temp_mem[4442];
   memory[1110][3] = temp_mem[4443];

   memory[1111][0] = temp_mem[4444];
   memory[1111][1] = temp_mem[4445];
   memory[1111][2] = temp_mem[4446];
   memory[1111][3] = temp_mem[4447];

   memory[1112][0] = temp_mem[4448];
   memory[1112][1] = temp_mem[4449];
   memory[1112][2] = temp_mem[4450];
   memory[1112][3] = temp_mem[4451];

   memory[1113][0] = temp_mem[4452];
   memory[1113][1] = temp_mem[4453];
   memory[1113][2] = temp_mem[4454];
   memory[1113][3] = temp_mem[4455];

   memory[1114][0] = temp_mem[4456];
   memory[1114][1] = temp_mem[4457];
   memory[1114][2] = temp_mem[4458];
   memory[1114][3] = temp_mem[4459];

   memory[1115][0] = temp_mem[4460];
   memory[1115][1] = temp_mem[4461];
   memory[1115][2] = temp_mem[4462];
   memory[1115][3] = temp_mem[4463];

   memory[1116][0] = temp_mem[4464];
   memory[1116][1] = temp_mem[4465];
   memory[1116][2] = temp_mem[4466];
   memory[1116][3] = temp_mem[4467];

   memory[1117][0] = temp_mem[4468];
   memory[1117][1] = temp_mem[4469];
   memory[1117][2] = temp_mem[4470];
   memory[1117][3] = temp_mem[4471];

   memory[1118][0] = temp_mem[4472];
   memory[1118][1] = temp_mem[4473];
   memory[1118][2] = temp_mem[4474];
   memory[1118][3] = temp_mem[4475];

   memory[1119][0] = temp_mem[4476];
   memory[1119][1] = temp_mem[4477];
   memory[1119][2] = temp_mem[4478];
   memory[1119][3] = temp_mem[4479];

   memory[1120][0] = temp_mem[4480];
   memory[1120][1] = temp_mem[4481];
   memory[1120][2] = temp_mem[4482];
   memory[1120][3] = temp_mem[4483];

   memory[1121][0] = temp_mem[4484];
   memory[1121][1] = temp_mem[4485];
   memory[1121][2] = temp_mem[4486];
   memory[1121][3] = temp_mem[4487];

   memory[1122][0] = temp_mem[4488];
   memory[1122][1] = temp_mem[4489];
   memory[1122][2] = temp_mem[4490];
   memory[1122][3] = temp_mem[4491];

   memory[1123][0] = temp_mem[4492];
   memory[1123][1] = temp_mem[4493];
   memory[1123][2] = temp_mem[4494];
   memory[1123][3] = temp_mem[4495];

   memory[1124][0] = temp_mem[4496];
   memory[1124][1] = temp_mem[4497];
   memory[1124][2] = temp_mem[4498];
   memory[1124][3] = temp_mem[4499];

   memory[1125][0] = temp_mem[4500];
   memory[1125][1] = temp_mem[4501];
   memory[1125][2] = temp_mem[4502];
   memory[1125][3] = temp_mem[4503];

   memory[1126][0] = temp_mem[4504];
   memory[1126][1] = temp_mem[4505];
   memory[1126][2] = temp_mem[4506];
   memory[1126][3] = temp_mem[4507];

   memory[1127][0] = temp_mem[4508];
   memory[1127][1] = temp_mem[4509];
   memory[1127][2] = temp_mem[4510];
   memory[1127][3] = temp_mem[4511];

   memory[1128][0] = temp_mem[4512];
   memory[1128][1] = temp_mem[4513];
   memory[1128][2] = temp_mem[4514];
   memory[1128][3] = temp_mem[4515];

   memory[1129][0] = temp_mem[4516];
   memory[1129][1] = temp_mem[4517];
   memory[1129][2] = temp_mem[4518];
   memory[1129][3] = temp_mem[4519];

   memory[1130][0] = temp_mem[4520];
   memory[1130][1] = temp_mem[4521];
   memory[1130][2] = temp_mem[4522];
   memory[1130][3] = temp_mem[4523];

   memory[1131][0] = temp_mem[4524];
   memory[1131][1] = temp_mem[4525];
   memory[1131][2] = temp_mem[4526];
   memory[1131][3] = temp_mem[4527];

   memory[1132][0] = temp_mem[4528];
   memory[1132][1] = temp_mem[4529];
   memory[1132][2] = temp_mem[4530];
   memory[1132][3] = temp_mem[4531];

   memory[1133][0] = temp_mem[4532];
   memory[1133][1] = temp_mem[4533];
   memory[1133][2] = temp_mem[4534];
   memory[1133][3] = temp_mem[4535];

   memory[1134][0] = temp_mem[4536];
   memory[1134][1] = temp_mem[4537];
   memory[1134][2] = temp_mem[4538];
   memory[1134][3] = temp_mem[4539];

   memory[1135][0] = temp_mem[4540];
   memory[1135][1] = temp_mem[4541];
   memory[1135][2] = temp_mem[4542];
   memory[1135][3] = temp_mem[4543];

   memory[1136][0] = temp_mem[4544];
   memory[1136][1] = temp_mem[4545];
   memory[1136][2] = temp_mem[4546];
   memory[1136][3] = temp_mem[4547];

   memory[1137][0] = temp_mem[4548];
   memory[1137][1] = temp_mem[4549];
   memory[1137][2] = temp_mem[4550];
   memory[1137][3] = temp_mem[4551];

   memory[1138][0] = temp_mem[4552];
   memory[1138][1] = temp_mem[4553];
   memory[1138][2] = temp_mem[4554];
   memory[1138][3] = temp_mem[4555];

   memory[1139][0] = temp_mem[4556];
   memory[1139][1] = temp_mem[4557];
   memory[1139][2] = temp_mem[4558];
   memory[1139][3] = temp_mem[4559];

   memory[1140][0] = temp_mem[4560];
   memory[1140][1] = temp_mem[4561];
   memory[1140][2] = temp_mem[4562];
   memory[1140][3] = temp_mem[4563];

   memory[1141][0] = temp_mem[4564];
   memory[1141][1] = temp_mem[4565];
   memory[1141][2] = temp_mem[4566];
   memory[1141][3] = temp_mem[4567];

   memory[1142][0] = temp_mem[4568];
   memory[1142][1] = temp_mem[4569];
   memory[1142][2] = temp_mem[4570];
   memory[1142][3] = temp_mem[4571];

   memory[1143][0] = temp_mem[4572];
   memory[1143][1] = temp_mem[4573];
   memory[1143][2] = temp_mem[4574];
   memory[1143][3] = temp_mem[4575];

   memory[1144][0] = temp_mem[4576];
   memory[1144][1] = temp_mem[4577];
   memory[1144][2] = temp_mem[4578];
   memory[1144][3] = temp_mem[4579];

   memory[1145][0] = temp_mem[4580];
   memory[1145][1] = temp_mem[4581];
   memory[1145][2] = temp_mem[4582];
   memory[1145][3] = temp_mem[4583];

   memory[1146][0] = temp_mem[4584];
   memory[1146][1] = temp_mem[4585];
   memory[1146][2] = temp_mem[4586];
   memory[1146][3] = temp_mem[4587];

   memory[1147][0] = temp_mem[4588];
   memory[1147][1] = temp_mem[4589];
   memory[1147][2] = temp_mem[4590];
   memory[1147][3] = temp_mem[4591];

   memory[1148][0] = temp_mem[4592];
   memory[1148][1] = temp_mem[4593];
   memory[1148][2] = temp_mem[4594];
   memory[1148][3] = temp_mem[4595];

   memory[1149][0] = temp_mem[4596];
   memory[1149][1] = temp_mem[4597];
   memory[1149][2] = temp_mem[4598];
   memory[1149][3] = temp_mem[4599];

   memory[1150][0] = temp_mem[4600];
   memory[1150][1] = temp_mem[4601];
   memory[1150][2] = temp_mem[4602];
   memory[1150][3] = temp_mem[4603];

   memory[1151][0] = temp_mem[4604];
   memory[1151][1] = temp_mem[4605];
   memory[1151][2] = temp_mem[4606];
   memory[1151][3] = temp_mem[4607];

   memory[1152][0] = temp_mem[4608];
   memory[1152][1] = temp_mem[4609];
   memory[1152][2] = temp_mem[4610];
   memory[1152][3] = temp_mem[4611];

   memory[1153][0] = temp_mem[4612];
   memory[1153][1] = temp_mem[4613];
   memory[1153][2] = temp_mem[4614];
   memory[1153][3] = temp_mem[4615];

   memory[1154][0] = temp_mem[4616];
   memory[1154][1] = temp_mem[4617];
   memory[1154][2] = temp_mem[4618];
   memory[1154][3] = temp_mem[4619];

   memory[1155][0] = temp_mem[4620];
   memory[1155][1] = temp_mem[4621];
   memory[1155][2] = temp_mem[4622];
   memory[1155][3] = temp_mem[4623];

   memory[1156][0] = temp_mem[4624];
   memory[1156][1] = temp_mem[4625];
   memory[1156][2] = temp_mem[4626];
   memory[1156][3] = temp_mem[4627];

   memory[1157][0] = temp_mem[4628];
   memory[1157][1] = temp_mem[4629];
   memory[1157][2] = temp_mem[4630];
   memory[1157][3] = temp_mem[4631];

   memory[1158][0] = temp_mem[4632];
   memory[1158][1] = temp_mem[4633];
   memory[1158][2] = temp_mem[4634];
   memory[1158][3] = temp_mem[4635];

   memory[1159][0] = temp_mem[4636];
   memory[1159][1] = temp_mem[4637];
   memory[1159][2] = temp_mem[4638];
   memory[1159][3] = temp_mem[4639];

   memory[1160][0] = temp_mem[4640];
   memory[1160][1] = temp_mem[4641];
   memory[1160][2] = temp_mem[4642];
   memory[1160][3] = temp_mem[4643];

   memory[1161][0] = temp_mem[4644];
   memory[1161][1] = temp_mem[4645];
   memory[1161][2] = temp_mem[4646];
   memory[1161][3] = temp_mem[4647];

   memory[1162][0] = temp_mem[4648];
   memory[1162][1] = temp_mem[4649];
   memory[1162][2] = temp_mem[4650];
   memory[1162][3] = temp_mem[4651];

   memory[1163][0] = temp_mem[4652];
   memory[1163][1] = temp_mem[4653];
   memory[1163][2] = temp_mem[4654];
   memory[1163][3] = temp_mem[4655];

   memory[1164][0] = temp_mem[4656];
   memory[1164][1] = temp_mem[4657];
   memory[1164][2] = temp_mem[4658];
   memory[1164][3] = temp_mem[4659];

   memory[1165][0] = temp_mem[4660];
   memory[1165][1] = temp_mem[4661];
   memory[1165][2] = temp_mem[4662];
   memory[1165][3] = temp_mem[4663];

   memory[1166][0] = temp_mem[4664];
   memory[1166][1] = temp_mem[4665];
   memory[1166][2] = temp_mem[4666];
   memory[1166][3] = temp_mem[4667];

   memory[1167][0] = temp_mem[4668];
   memory[1167][1] = temp_mem[4669];
   memory[1167][2] = temp_mem[4670];
   memory[1167][3] = temp_mem[4671];

   memory[1168][0] = temp_mem[4672];
   memory[1168][1] = temp_mem[4673];
   memory[1168][2] = temp_mem[4674];
   memory[1168][3] = temp_mem[4675];

   memory[1169][0] = temp_mem[4676];
   memory[1169][1] = temp_mem[4677];
   memory[1169][2] = temp_mem[4678];
   memory[1169][3] = temp_mem[4679];

   memory[1170][0] = temp_mem[4680];
   memory[1170][1] = temp_mem[4681];
   memory[1170][2] = temp_mem[4682];
   memory[1170][3] = temp_mem[4683];

   memory[1171][0] = temp_mem[4684];
   memory[1171][1] = temp_mem[4685];
   memory[1171][2] = temp_mem[4686];
   memory[1171][3] = temp_mem[4687];

   memory[1172][0] = temp_mem[4688];
   memory[1172][1] = temp_mem[4689];
   memory[1172][2] = temp_mem[4690];
   memory[1172][3] = temp_mem[4691];

   memory[1173][0] = temp_mem[4692];
   memory[1173][1] = temp_mem[4693];
   memory[1173][2] = temp_mem[4694];
   memory[1173][3] = temp_mem[4695];

   memory[1174][0] = temp_mem[4696];
   memory[1174][1] = temp_mem[4697];
   memory[1174][2] = temp_mem[4698];
   memory[1174][3] = temp_mem[4699];

   memory[1175][0] = temp_mem[4700];
   memory[1175][1] = temp_mem[4701];
   memory[1175][2] = temp_mem[4702];
   memory[1175][3] = temp_mem[4703];

   memory[1176][0] = temp_mem[4704];
   memory[1176][1] = temp_mem[4705];
   memory[1176][2] = temp_mem[4706];
   memory[1176][3] = temp_mem[4707];

   memory[1177][0] = temp_mem[4708];
   memory[1177][1] = temp_mem[4709];
   memory[1177][2] = temp_mem[4710];
   memory[1177][3] = temp_mem[4711];

   memory[1178][0] = temp_mem[4712];
   memory[1178][1] = temp_mem[4713];
   memory[1178][2] = temp_mem[4714];
   memory[1178][3] = temp_mem[4715];

   memory[1179][0] = temp_mem[4716];
   memory[1179][1] = temp_mem[4717];
   memory[1179][2] = temp_mem[4718];
   memory[1179][3] = temp_mem[4719];

   memory[1180][0] = temp_mem[4720];
   memory[1180][1] = temp_mem[4721];
   memory[1180][2] = temp_mem[4722];
   memory[1180][3] = temp_mem[4723];

   memory[1181][0] = temp_mem[4724];
   memory[1181][1] = temp_mem[4725];
   memory[1181][2] = temp_mem[4726];
   memory[1181][3] = temp_mem[4727];

   memory[1182][0] = temp_mem[4728];
   memory[1182][1] = temp_mem[4729];
   memory[1182][2] = temp_mem[4730];
   memory[1182][3] = temp_mem[4731];

   memory[1183][0] = temp_mem[4732];
   memory[1183][1] = temp_mem[4733];
   memory[1183][2] = temp_mem[4734];
   memory[1183][3] = temp_mem[4735];

   memory[1184][0] = temp_mem[4736];
   memory[1184][1] = temp_mem[4737];
   memory[1184][2] = temp_mem[4738];
   memory[1184][3] = temp_mem[4739];

   memory[1185][0] = temp_mem[4740];
   memory[1185][1] = temp_mem[4741];
   memory[1185][2] = temp_mem[4742];
   memory[1185][3] = temp_mem[4743];

   memory[1186][0] = temp_mem[4744];
   memory[1186][1] = temp_mem[4745];
   memory[1186][2] = temp_mem[4746];
   memory[1186][3] = temp_mem[4747];

   memory[1187][0] = temp_mem[4748];
   memory[1187][1] = temp_mem[4749];
   memory[1187][2] = temp_mem[4750];
   memory[1187][3] = temp_mem[4751];

   memory[1188][0] = temp_mem[4752];
   memory[1188][1] = temp_mem[4753];
   memory[1188][2] = temp_mem[4754];
   memory[1188][3] = temp_mem[4755];

   memory[1189][0] = temp_mem[4756];
   memory[1189][1] = temp_mem[4757];
   memory[1189][2] = temp_mem[4758];
   memory[1189][3] = temp_mem[4759];

   memory[1190][0] = temp_mem[4760];
   memory[1190][1] = temp_mem[4761];
   memory[1190][2] = temp_mem[4762];
   memory[1190][3] = temp_mem[4763];

   memory[1191][0] = temp_mem[4764];
   memory[1191][1] = temp_mem[4765];
   memory[1191][2] = temp_mem[4766];
   memory[1191][3] = temp_mem[4767];

   memory[1192][0] = temp_mem[4768];
   memory[1192][1] = temp_mem[4769];
   memory[1192][2] = temp_mem[4770];
   memory[1192][3] = temp_mem[4771];

   memory[1193][0] = temp_mem[4772];
   memory[1193][1] = temp_mem[4773];
   memory[1193][2] = temp_mem[4774];
   memory[1193][3] = temp_mem[4775];

   memory[1194][0] = temp_mem[4776];
   memory[1194][1] = temp_mem[4777];
   memory[1194][2] = temp_mem[4778];
   memory[1194][3] = temp_mem[4779];

   memory[1195][0] = temp_mem[4780];
   memory[1195][1] = temp_mem[4781];
   memory[1195][2] = temp_mem[4782];
   memory[1195][3] = temp_mem[4783];

   memory[1196][0] = temp_mem[4784];
   memory[1196][1] = temp_mem[4785];
   memory[1196][2] = temp_mem[4786];
   memory[1196][3] = temp_mem[4787];

   memory[1197][0] = temp_mem[4788];
   memory[1197][1] = temp_mem[4789];
   memory[1197][2] = temp_mem[4790];
   memory[1197][3] = temp_mem[4791];

   memory[1198][0] = temp_mem[4792];
   memory[1198][1] = temp_mem[4793];
   memory[1198][2] = temp_mem[4794];
   memory[1198][3] = temp_mem[4795];

   memory[1199][0] = temp_mem[4796];
   memory[1199][1] = temp_mem[4797];
   memory[1199][2] = temp_mem[4798];
   memory[1199][3] = temp_mem[4799];

   memory[1200][0] = temp_mem[4800];
   memory[1200][1] = temp_mem[4801];
   memory[1200][2] = temp_mem[4802];
   memory[1200][3] = temp_mem[4803];

   memory[1201][0] = temp_mem[4804];
   memory[1201][1] = temp_mem[4805];
   memory[1201][2] = temp_mem[4806];
   memory[1201][3] = temp_mem[4807];

   memory[1202][0] = temp_mem[4808];
   memory[1202][1] = temp_mem[4809];
   memory[1202][2] = temp_mem[4810];
   memory[1202][3] = temp_mem[4811];

   memory[1203][0] = temp_mem[4812];
   memory[1203][1] = temp_mem[4813];
   memory[1203][2] = temp_mem[4814];
   memory[1203][3] = temp_mem[4815];

   memory[1204][0] = temp_mem[4816];
   memory[1204][1] = temp_mem[4817];
   memory[1204][2] = temp_mem[4818];
   memory[1204][3] = temp_mem[4819];

   memory[1205][0] = temp_mem[4820];
   memory[1205][1] = temp_mem[4821];
   memory[1205][2] = temp_mem[4822];
   memory[1205][3] = temp_mem[4823];

   memory[1206][0] = temp_mem[4824];
   memory[1206][1] = temp_mem[4825];
   memory[1206][2] = temp_mem[4826];
   memory[1206][3] = temp_mem[4827];

   memory[1207][0] = temp_mem[4828];
   memory[1207][1] = temp_mem[4829];
   memory[1207][2] = temp_mem[4830];
   memory[1207][3] = temp_mem[4831];

   memory[1208][0] = temp_mem[4832];
   memory[1208][1] = temp_mem[4833];
   memory[1208][2] = temp_mem[4834];
   memory[1208][3] = temp_mem[4835];

   memory[1209][0] = temp_mem[4836];
   memory[1209][1] = temp_mem[4837];
   memory[1209][2] = temp_mem[4838];
   memory[1209][3] = temp_mem[4839];

   memory[1210][0] = temp_mem[4840];
   memory[1210][1] = temp_mem[4841];
   memory[1210][2] = temp_mem[4842];
   memory[1210][3] = temp_mem[4843];

   memory[1211][0] = temp_mem[4844];
   memory[1211][1] = temp_mem[4845];
   memory[1211][2] = temp_mem[4846];
   memory[1211][3] = temp_mem[4847];

   memory[1212][0] = temp_mem[4848];
   memory[1212][1] = temp_mem[4849];
   memory[1212][2] = temp_mem[4850];
   memory[1212][3] = temp_mem[4851];

   memory[1213][0] = temp_mem[4852];
   memory[1213][1] = temp_mem[4853];
   memory[1213][2] = temp_mem[4854];
   memory[1213][3] = temp_mem[4855];

   memory[1214][0] = temp_mem[4856];
   memory[1214][1] = temp_mem[4857];
   memory[1214][2] = temp_mem[4858];
   memory[1214][3] = temp_mem[4859];

   memory[1215][0] = temp_mem[4860];
   memory[1215][1] = temp_mem[4861];
   memory[1215][2] = temp_mem[4862];
   memory[1215][3] = temp_mem[4863];

   memory[1216][0] = temp_mem[4864];
   memory[1216][1] = temp_mem[4865];
   memory[1216][2] = temp_mem[4866];
   memory[1216][3] = temp_mem[4867];

   memory[1217][0] = temp_mem[4868];
   memory[1217][1] = temp_mem[4869];
   memory[1217][2] = temp_mem[4870];
   memory[1217][3] = temp_mem[4871];

   memory[1218][0] = temp_mem[4872];
   memory[1218][1] = temp_mem[4873];
   memory[1218][2] = temp_mem[4874];
   memory[1218][3] = temp_mem[4875];

   memory[1219][0] = temp_mem[4876];
   memory[1219][1] = temp_mem[4877];
   memory[1219][2] = temp_mem[4878];
   memory[1219][3] = temp_mem[4879];

   memory[1220][0] = temp_mem[4880];
   memory[1220][1] = temp_mem[4881];
   memory[1220][2] = temp_mem[4882];
   memory[1220][3] = temp_mem[4883];

   memory[1221][0] = temp_mem[4884];
   memory[1221][1] = temp_mem[4885];
   memory[1221][2] = temp_mem[4886];
   memory[1221][3] = temp_mem[4887];

   memory[1222][0] = temp_mem[4888];
   memory[1222][1] = temp_mem[4889];
   memory[1222][2] = temp_mem[4890];
   memory[1222][3] = temp_mem[4891];

   memory[1223][0] = temp_mem[4892];
   memory[1223][1] = temp_mem[4893];
   memory[1223][2] = temp_mem[4894];
   memory[1223][3] = temp_mem[4895];

   memory[1224][0] = temp_mem[4896];
   memory[1224][1] = temp_mem[4897];
   memory[1224][2] = temp_mem[4898];
   memory[1224][3] = temp_mem[4899];

   memory[1225][0] = temp_mem[4900];
   memory[1225][1] = temp_mem[4901];
   memory[1225][2] = temp_mem[4902];
   memory[1225][3] = temp_mem[4903];

   memory[1226][0] = temp_mem[4904];
   memory[1226][1] = temp_mem[4905];
   memory[1226][2] = temp_mem[4906];
   memory[1226][3] = temp_mem[4907];

   memory[1227][0] = temp_mem[4908];
   memory[1227][1] = temp_mem[4909];
   memory[1227][2] = temp_mem[4910];
   memory[1227][3] = temp_mem[4911];

   memory[1228][0] = temp_mem[4912];
   memory[1228][1] = temp_mem[4913];
   memory[1228][2] = temp_mem[4914];
   memory[1228][3] = temp_mem[4915];

   memory[1229][0] = temp_mem[4916];
   memory[1229][1] = temp_mem[4917];
   memory[1229][2] = temp_mem[4918];
   memory[1229][3] = temp_mem[4919];

   memory[1230][0] = temp_mem[4920];
   memory[1230][1] = temp_mem[4921];
   memory[1230][2] = temp_mem[4922];
   memory[1230][3] = temp_mem[4923];

   memory[1231][0] = temp_mem[4924];
   memory[1231][1] = temp_mem[4925];
   memory[1231][2] = temp_mem[4926];
   memory[1231][3] = temp_mem[4927];

   memory[1232][0] = temp_mem[4928];
   memory[1232][1] = temp_mem[4929];
   memory[1232][2] = temp_mem[4930];
   memory[1232][3] = temp_mem[4931];

   memory[1233][0] = temp_mem[4932];
   memory[1233][1] = temp_mem[4933];
   memory[1233][2] = temp_mem[4934];
   memory[1233][3] = temp_mem[4935];

   memory[1234][0] = temp_mem[4936];
   memory[1234][1] = temp_mem[4937];
   memory[1234][2] = temp_mem[4938];
   memory[1234][3] = temp_mem[4939];

   memory[1235][0] = temp_mem[4940];
   memory[1235][1] = temp_mem[4941];
   memory[1235][2] = temp_mem[4942];
   memory[1235][3] = temp_mem[4943];

   memory[1236][0] = temp_mem[4944];
   memory[1236][1] = temp_mem[4945];
   memory[1236][2] = temp_mem[4946];
   memory[1236][3] = temp_mem[4947];

   memory[1237][0] = temp_mem[4948];
   memory[1237][1] = temp_mem[4949];
   memory[1237][2] = temp_mem[4950];
   memory[1237][3] = temp_mem[4951];

   memory[1238][0] = temp_mem[4952];
   memory[1238][1] = temp_mem[4953];
   memory[1238][2] = temp_mem[4954];
   memory[1238][3] = temp_mem[4955];

   memory[1239][0] = temp_mem[4956];
   memory[1239][1] = temp_mem[4957];
   memory[1239][2] = temp_mem[4958];
   memory[1239][3] = temp_mem[4959];

   memory[1240][0] = temp_mem[4960];
   memory[1240][1] = temp_mem[4961];
   memory[1240][2] = temp_mem[4962];
   memory[1240][3] = temp_mem[4963];

   memory[1241][0] = temp_mem[4964];
   memory[1241][1] = temp_mem[4965];
   memory[1241][2] = temp_mem[4966];
   memory[1241][3] = temp_mem[4967];

   memory[1242][0] = temp_mem[4968];
   memory[1242][1] = temp_mem[4969];
   memory[1242][2] = temp_mem[4970];
   memory[1242][3] = temp_mem[4971];

   memory[1243][0] = temp_mem[4972];
   memory[1243][1] = temp_mem[4973];
   memory[1243][2] = temp_mem[4974];
   memory[1243][3] = temp_mem[4975];

   memory[1244][0] = temp_mem[4976];
   memory[1244][1] = temp_mem[4977];
   memory[1244][2] = temp_mem[4978];
   memory[1244][3] = temp_mem[4979];

   memory[1245][0] = temp_mem[4980];
   memory[1245][1] = temp_mem[4981];
   memory[1245][2] = temp_mem[4982];
   memory[1245][3] = temp_mem[4983];

   memory[1246][0] = temp_mem[4984];
   memory[1246][1] = temp_mem[4985];
   memory[1246][2] = temp_mem[4986];
   memory[1246][3] = temp_mem[4987];

   memory[1247][0] = temp_mem[4988];
   memory[1247][1] = temp_mem[4989];
   memory[1247][2] = temp_mem[4990];
   memory[1247][3] = temp_mem[4991];

   memory[1248][0] = temp_mem[4992];
   memory[1248][1] = temp_mem[4993];
   memory[1248][2] = temp_mem[4994];
   memory[1248][3] = temp_mem[4995];

   memory[1249][0] = temp_mem[4996];
   memory[1249][1] = temp_mem[4997];
   memory[1249][2] = temp_mem[4998];
   memory[1249][3] = temp_mem[4999];

   memory[1250][0] = temp_mem[5000];
   memory[1250][1] = temp_mem[5001];
   memory[1250][2] = temp_mem[5002];
   memory[1250][3] = temp_mem[5003];

   memory[1251][0] = temp_mem[5004];
   memory[1251][1] = temp_mem[5005];
   memory[1251][2] = temp_mem[5006];
   memory[1251][3] = temp_mem[5007];

   memory[1252][0] = temp_mem[5008];
   memory[1252][1] = temp_mem[5009];
   memory[1252][2] = temp_mem[5010];
   memory[1252][3] = temp_mem[5011];

   memory[1253][0] = temp_mem[5012];
   memory[1253][1] = temp_mem[5013];
   memory[1253][2] = temp_mem[5014];
   memory[1253][3] = temp_mem[5015];

   memory[1254][0] = temp_mem[5016];
   memory[1254][1] = temp_mem[5017];
   memory[1254][2] = temp_mem[5018];
   memory[1254][3] = temp_mem[5019];

   memory[1255][0] = temp_mem[5020];
   memory[1255][1] = temp_mem[5021];
   memory[1255][2] = temp_mem[5022];
   memory[1255][3] = temp_mem[5023];

   memory[1256][0] = temp_mem[5024];
   memory[1256][1] = temp_mem[5025];
   memory[1256][2] = temp_mem[5026];
   memory[1256][3] = temp_mem[5027];

   memory[1257][0] = temp_mem[5028];
   memory[1257][1] = temp_mem[5029];
   memory[1257][2] = temp_mem[5030];
   memory[1257][3] = temp_mem[5031];

   memory[1258][0] = temp_mem[5032];
   memory[1258][1] = temp_mem[5033];
   memory[1258][2] = temp_mem[5034];
   memory[1258][3] = temp_mem[5035];

   memory[1259][0] = temp_mem[5036];
   memory[1259][1] = temp_mem[5037];
   memory[1259][2] = temp_mem[5038];
   memory[1259][3] = temp_mem[5039];

   memory[1260][0] = temp_mem[5040];
   memory[1260][1] = temp_mem[5041];
   memory[1260][2] = temp_mem[5042];
   memory[1260][3] = temp_mem[5043];

   memory[1261][0] = temp_mem[5044];
   memory[1261][1] = temp_mem[5045];
   memory[1261][2] = temp_mem[5046];
   memory[1261][3] = temp_mem[5047];

   memory[1262][0] = temp_mem[5048];
   memory[1262][1] = temp_mem[5049];
   memory[1262][2] = temp_mem[5050];
   memory[1262][3] = temp_mem[5051];

   memory[1263][0] = temp_mem[5052];
   memory[1263][1] = temp_mem[5053];
   memory[1263][2] = temp_mem[5054];
   memory[1263][3] = temp_mem[5055];

   memory[1264][0] = temp_mem[5056];
   memory[1264][1] = temp_mem[5057];
   memory[1264][2] = temp_mem[5058];
   memory[1264][3] = temp_mem[5059];

   memory[1265][0] = temp_mem[5060];
   memory[1265][1] = temp_mem[5061];
   memory[1265][2] = temp_mem[5062];
   memory[1265][3] = temp_mem[5063];

   memory[1266][0] = temp_mem[5064];
   memory[1266][1] = temp_mem[5065];
   memory[1266][2] = temp_mem[5066];
   memory[1266][3] = temp_mem[5067];

   memory[1267][0] = temp_mem[5068];
   memory[1267][1] = temp_mem[5069];
   memory[1267][2] = temp_mem[5070];
   memory[1267][3] = temp_mem[5071];

   memory[1268][0] = temp_mem[5072];
   memory[1268][1] = temp_mem[5073];
   memory[1268][2] = temp_mem[5074];
   memory[1268][3] = temp_mem[5075];

   memory[1269][0] = temp_mem[5076];
   memory[1269][1] = temp_mem[5077];
   memory[1269][2] = temp_mem[5078];
   memory[1269][3] = temp_mem[5079];

   memory[1270][0] = temp_mem[5080];
   memory[1270][1] = temp_mem[5081];
   memory[1270][2] = temp_mem[5082];
   memory[1270][3] = temp_mem[5083];

   memory[1271][0] = temp_mem[5084];
   memory[1271][1] = temp_mem[5085];
   memory[1271][2] = temp_mem[5086];
   memory[1271][3] = temp_mem[5087];

   memory[1272][0] = temp_mem[5088];
   memory[1272][1] = temp_mem[5089];
   memory[1272][2] = temp_mem[5090];
   memory[1272][3] = temp_mem[5091];

   memory[1273][0] = temp_mem[5092];
   memory[1273][1] = temp_mem[5093];
   memory[1273][2] = temp_mem[5094];
   memory[1273][3] = temp_mem[5095];

   memory[1274][0] = temp_mem[5096];
   memory[1274][1] = temp_mem[5097];
   memory[1274][2] = temp_mem[5098];
   memory[1274][3] = temp_mem[5099];

   memory[1275][0] = temp_mem[5100];
   memory[1275][1] = temp_mem[5101];
   memory[1275][2] = temp_mem[5102];
   memory[1275][3] = temp_mem[5103];

   memory[1276][0] = temp_mem[5104];
   memory[1276][1] = temp_mem[5105];
   memory[1276][2] = temp_mem[5106];
   memory[1276][3] = temp_mem[5107];

   memory[1277][0] = temp_mem[5108];
   memory[1277][1] = temp_mem[5109];
   memory[1277][2] = temp_mem[5110];
   memory[1277][3] = temp_mem[5111];

   memory[1278][0] = temp_mem[5112];
   memory[1278][1] = temp_mem[5113];
   memory[1278][2] = temp_mem[5114];
   memory[1278][3] = temp_mem[5115];

   memory[1279][0] = temp_mem[5116];
   memory[1279][1] = temp_mem[5117];
   memory[1279][2] = temp_mem[5118];
   memory[1279][3] = temp_mem[5119];

   memory[1280][0] = temp_mem[5120];
   memory[1280][1] = temp_mem[5121];
   memory[1280][2] = temp_mem[5122];
   memory[1280][3] = temp_mem[5123];

   memory[1281][0] = temp_mem[5124];
   memory[1281][1] = temp_mem[5125];
   memory[1281][2] = temp_mem[5126];
   memory[1281][3] = temp_mem[5127];

   memory[1282][0] = temp_mem[5128];
   memory[1282][1] = temp_mem[5129];
   memory[1282][2] = temp_mem[5130];
   memory[1282][3] = temp_mem[5131];

   memory[1283][0] = temp_mem[5132];
   memory[1283][1] = temp_mem[5133];
   memory[1283][2] = temp_mem[5134];
   memory[1283][3] = temp_mem[5135];

   memory[1284][0] = temp_mem[5136];
   memory[1284][1] = temp_mem[5137];
   memory[1284][2] = temp_mem[5138];
   memory[1284][3] = temp_mem[5139];

   memory[1285][0] = temp_mem[5140];
   memory[1285][1] = temp_mem[5141];
   memory[1285][2] = temp_mem[5142];
   memory[1285][3] = temp_mem[5143];

   memory[1286][0] = temp_mem[5144];
   memory[1286][1] = temp_mem[5145];
   memory[1286][2] = temp_mem[5146];
   memory[1286][3] = temp_mem[5147];

   memory[1287][0] = temp_mem[5148];
   memory[1287][1] = temp_mem[5149];
   memory[1287][2] = temp_mem[5150];
   memory[1287][3] = temp_mem[5151];

   memory[1288][0] = temp_mem[5152];
   memory[1288][1] = temp_mem[5153];
   memory[1288][2] = temp_mem[5154];
   memory[1288][3] = temp_mem[5155];

   memory[1289][0] = temp_mem[5156];
   memory[1289][1] = temp_mem[5157];
   memory[1289][2] = temp_mem[5158];
   memory[1289][3] = temp_mem[5159];

   memory[1290][0] = temp_mem[5160];
   memory[1290][1] = temp_mem[5161];
   memory[1290][2] = temp_mem[5162];
   memory[1290][3] = temp_mem[5163];

   memory[1291][0] = temp_mem[5164];
   memory[1291][1] = temp_mem[5165];
   memory[1291][2] = temp_mem[5166];
   memory[1291][3] = temp_mem[5167];

   memory[1292][0] = temp_mem[5168];
   memory[1292][1] = temp_mem[5169];
   memory[1292][2] = temp_mem[5170];
   memory[1292][3] = temp_mem[5171];

   memory[1293][0] = temp_mem[5172];
   memory[1293][1] = temp_mem[5173];
   memory[1293][2] = temp_mem[5174];
   memory[1293][3] = temp_mem[5175];

   memory[1294][0] = temp_mem[5176];
   memory[1294][1] = temp_mem[5177];
   memory[1294][2] = temp_mem[5178];
   memory[1294][3] = temp_mem[5179];

   memory[1295][0] = temp_mem[5180];
   memory[1295][1] = temp_mem[5181];
   memory[1295][2] = temp_mem[5182];
   memory[1295][3] = temp_mem[5183];

   memory[1296][0] = temp_mem[5184];
   memory[1296][1] = temp_mem[5185];
   memory[1296][2] = temp_mem[5186];
   memory[1296][3] = temp_mem[5187];

   memory[1297][0] = temp_mem[5188];
   memory[1297][1] = temp_mem[5189];
   memory[1297][2] = temp_mem[5190];
   memory[1297][3] = temp_mem[5191];

   memory[1298][0] = temp_mem[5192];
   memory[1298][1] = temp_mem[5193];
   memory[1298][2] = temp_mem[5194];
   memory[1298][3] = temp_mem[5195];

   memory[1299][0] = temp_mem[5196];
   memory[1299][1] = temp_mem[5197];
   memory[1299][2] = temp_mem[5198];
   memory[1299][3] = temp_mem[5199];

   memory[1300][0] = temp_mem[5200];
   memory[1300][1] = temp_mem[5201];
   memory[1300][2] = temp_mem[5202];
   memory[1300][3] = temp_mem[5203];

   memory[1301][0] = temp_mem[5204];
   memory[1301][1] = temp_mem[5205];
   memory[1301][2] = temp_mem[5206];
   memory[1301][3] = temp_mem[5207];

   memory[1302][0] = temp_mem[5208];
   memory[1302][1] = temp_mem[5209];
   memory[1302][2] = temp_mem[5210];
   memory[1302][3] = temp_mem[5211];

   memory[1303][0] = temp_mem[5212];
   memory[1303][1] = temp_mem[5213];
   memory[1303][2] = temp_mem[5214];
   memory[1303][3] = temp_mem[5215];

   memory[1304][0] = temp_mem[5216];
   memory[1304][1] = temp_mem[5217];
   memory[1304][2] = temp_mem[5218];
   memory[1304][3] = temp_mem[5219];

   memory[1305][0] = temp_mem[5220];
   memory[1305][1] = temp_mem[5221];
   memory[1305][2] = temp_mem[5222];
   memory[1305][3] = temp_mem[5223];

   memory[1306][0] = temp_mem[5224];
   memory[1306][1] = temp_mem[5225];
   memory[1306][2] = temp_mem[5226];
   memory[1306][3] = temp_mem[5227];

   memory[1307][0] = temp_mem[5228];
   memory[1307][1] = temp_mem[5229];
   memory[1307][2] = temp_mem[5230];
   memory[1307][3] = temp_mem[5231];

   memory[1308][0] = temp_mem[5232];
   memory[1308][1] = temp_mem[5233];
   memory[1308][2] = temp_mem[5234];
   memory[1308][3] = temp_mem[5235];

   memory[1309][0] = temp_mem[5236];
   memory[1309][1] = temp_mem[5237];
   memory[1309][2] = temp_mem[5238];
   memory[1309][3] = temp_mem[5239];

   memory[1310][0] = temp_mem[5240];
   memory[1310][1] = temp_mem[5241];
   memory[1310][2] = temp_mem[5242];
   memory[1310][3] = temp_mem[5243];

   memory[1311][0] = temp_mem[5244];
   memory[1311][1] = temp_mem[5245];
   memory[1311][2] = temp_mem[5246];
   memory[1311][3] = temp_mem[5247];

   memory[1312][0] = temp_mem[5248];
   memory[1312][1] = temp_mem[5249];
   memory[1312][2] = temp_mem[5250];
   memory[1312][3] = temp_mem[5251];

   memory[1313][0] = temp_mem[5252];
   memory[1313][1] = temp_mem[5253];
   memory[1313][2] = temp_mem[5254];
   memory[1313][3] = temp_mem[5255];

   memory[1314][0] = temp_mem[5256];
   memory[1314][1] = temp_mem[5257];
   memory[1314][2] = temp_mem[5258];
   memory[1314][3] = temp_mem[5259];

   memory[1315][0] = temp_mem[5260];
   memory[1315][1] = temp_mem[5261];
   memory[1315][2] = temp_mem[5262];
   memory[1315][3] = temp_mem[5263];

   memory[1316][0] = temp_mem[5264];
   memory[1316][1] = temp_mem[5265];
   memory[1316][2] = temp_mem[5266];
   memory[1316][3] = temp_mem[5267];

   memory[1317][0] = temp_mem[5268];
   memory[1317][1] = temp_mem[5269];
   memory[1317][2] = temp_mem[5270];
   memory[1317][3] = temp_mem[5271];

   memory[1318][0] = temp_mem[5272];
   memory[1318][1] = temp_mem[5273];
   memory[1318][2] = temp_mem[5274];
   memory[1318][3] = temp_mem[5275];

   memory[1319][0] = temp_mem[5276];
   memory[1319][1] = temp_mem[5277];
   memory[1319][2] = temp_mem[5278];
   memory[1319][3] = temp_mem[5279];

   memory[1320][0] = temp_mem[5280];
   memory[1320][1] = temp_mem[5281];
   memory[1320][2] = temp_mem[5282];
   memory[1320][3] = temp_mem[5283];

   memory[1321][0] = temp_mem[5284];
   memory[1321][1] = temp_mem[5285];
   memory[1321][2] = temp_mem[5286];
   memory[1321][3] = temp_mem[5287];

   memory[1322][0] = temp_mem[5288];
   memory[1322][1] = temp_mem[5289];
   memory[1322][2] = temp_mem[5290];
   memory[1322][3] = temp_mem[5291];

   memory[1323][0] = temp_mem[5292];
   memory[1323][1] = temp_mem[5293];
   memory[1323][2] = temp_mem[5294];
   memory[1323][3] = temp_mem[5295];

   memory[1324][0] = temp_mem[5296];
   memory[1324][1] = temp_mem[5297];
   memory[1324][2] = temp_mem[5298];
   memory[1324][3] = temp_mem[5299];

   memory[1325][0] = temp_mem[5300];
   memory[1325][1] = temp_mem[5301];
   memory[1325][2] = temp_mem[5302];
   memory[1325][3] = temp_mem[5303];

   memory[1326][0] = temp_mem[5304];
   memory[1326][1] = temp_mem[5305];
   memory[1326][2] = temp_mem[5306];
   memory[1326][3] = temp_mem[5307];

   memory[1327][0] = temp_mem[5308];
   memory[1327][1] = temp_mem[5309];
   memory[1327][2] = temp_mem[5310];
   memory[1327][3] = temp_mem[5311];

   memory[1328][0] = temp_mem[5312];
   memory[1328][1] = temp_mem[5313];
   memory[1328][2] = temp_mem[5314];
   memory[1328][3] = temp_mem[5315];

   memory[1329][0] = temp_mem[5316];
   memory[1329][1] = temp_mem[5317];
   memory[1329][2] = temp_mem[5318];
   memory[1329][3] = temp_mem[5319];

   memory[1330][0] = temp_mem[5320];
   memory[1330][1] = temp_mem[5321];
   memory[1330][2] = temp_mem[5322];
   memory[1330][3] = temp_mem[5323];

   memory[1331][0] = temp_mem[5324];
   memory[1331][1] = temp_mem[5325];
   memory[1331][2] = temp_mem[5326];
   memory[1331][3] = temp_mem[5327];

   memory[1332][0] = temp_mem[5328];
   memory[1332][1] = temp_mem[5329];
   memory[1332][2] = temp_mem[5330];
   memory[1332][3] = temp_mem[5331];

   memory[1333][0] = temp_mem[5332];
   memory[1333][1] = temp_mem[5333];
   memory[1333][2] = temp_mem[5334];
   memory[1333][3] = temp_mem[5335];

   memory[1334][0] = temp_mem[5336];
   memory[1334][1] = temp_mem[5337];
   memory[1334][2] = temp_mem[5338];
   memory[1334][3] = temp_mem[5339];

   memory[1335][0] = temp_mem[5340];
   memory[1335][1] = temp_mem[5341];
   memory[1335][2] = temp_mem[5342];
   memory[1335][3] = temp_mem[5343];

   memory[1336][0] = temp_mem[5344];
   memory[1336][1] = temp_mem[5345];
   memory[1336][2] = temp_mem[5346];
   memory[1336][3] = temp_mem[5347];

   memory[1337][0] = temp_mem[5348];
   memory[1337][1] = temp_mem[5349];
   memory[1337][2] = temp_mem[5350];
   memory[1337][3] = temp_mem[5351];

   memory[1338][0] = temp_mem[5352];
   memory[1338][1] = temp_mem[5353];
   memory[1338][2] = temp_mem[5354];
   memory[1338][3] = temp_mem[5355];

   memory[1339][0] = temp_mem[5356];
   memory[1339][1] = temp_mem[5357];
   memory[1339][2] = temp_mem[5358];
   memory[1339][3] = temp_mem[5359];

   memory[1340][0] = temp_mem[5360];
   memory[1340][1] = temp_mem[5361];
   memory[1340][2] = temp_mem[5362];
   memory[1340][3] = temp_mem[5363];

   memory[1341][0] = temp_mem[5364];
   memory[1341][1] = temp_mem[5365];
   memory[1341][2] = temp_mem[5366];
   memory[1341][3] = temp_mem[5367];

   memory[1342][0] = temp_mem[5368];
   memory[1342][1] = temp_mem[5369];
   memory[1342][2] = temp_mem[5370];
   memory[1342][3] = temp_mem[5371];

   memory[1343][0] = temp_mem[5372];
   memory[1343][1] = temp_mem[5373];
   memory[1343][2] = temp_mem[5374];
   memory[1343][3] = temp_mem[5375];

   memory[1344][0] = temp_mem[5376];
   memory[1344][1] = temp_mem[5377];
   memory[1344][2] = temp_mem[5378];
   memory[1344][3] = temp_mem[5379];

   memory[1345][0] = temp_mem[5380];
   memory[1345][1] = temp_mem[5381];
   memory[1345][2] = temp_mem[5382];
   memory[1345][3] = temp_mem[5383];

   memory[1346][0] = temp_mem[5384];
   memory[1346][1] = temp_mem[5385];
   memory[1346][2] = temp_mem[5386];
   memory[1346][3] = temp_mem[5387];

   memory[1347][0] = temp_mem[5388];
   memory[1347][1] = temp_mem[5389];
   memory[1347][2] = temp_mem[5390];
   memory[1347][3] = temp_mem[5391];

   memory[1348][0] = temp_mem[5392];
   memory[1348][1] = temp_mem[5393];
   memory[1348][2] = temp_mem[5394];
   memory[1348][3] = temp_mem[5395];

   memory[1349][0] = temp_mem[5396];
   memory[1349][1] = temp_mem[5397];
   memory[1349][2] = temp_mem[5398];
   memory[1349][3] = temp_mem[5399];

   memory[1350][0] = temp_mem[5400];
   memory[1350][1] = temp_mem[5401];
   memory[1350][2] = temp_mem[5402];
   memory[1350][3] = temp_mem[5403];

   memory[1351][0] = temp_mem[5404];
   memory[1351][1] = temp_mem[5405];
   memory[1351][2] = temp_mem[5406];
   memory[1351][3] = temp_mem[5407];

   memory[1352][0] = temp_mem[5408];
   memory[1352][1] = temp_mem[5409];
   memory[1352][2] = temp_mem[5410];
   memory[1352][3] = temp_mem[5411];

   memory[1353][0] = temp_mem[5412];
   memory[1353][1] = temp_mem[5413];
   memory[1353][2] = temp_mem[5414];
   memory[1353][3] = temp_mem[5415];

   memory[1354][0] = temp_mem[5416];
   memory[1354][1] = temp_mem[5417];
   memory[1354][2] = temp_mem[5418];
   memory[1354][3] = temp_mem[5419];

   memory[1355][0] = temp_mem[5420];
   memory[1355][1] = temp_mem[5421];
   memory[1355][2] = temp_mem[5422];
   memory[1355][3] = temp_mem[5423];

   memory[1356][0] = temp_mem[5424];
   memory[1356][1] = temp_mem[5425];
   memory[1356][2] = temp_mem[5426];
   memory[1356][3] = temp_mem[5427];

   memory[1357][0] = temp_mem[5428];
   memory[1357][1] = temp_mem[5429];
   memory[1357][2] = temp_mem[5430];
   memory[1357][3] = temp_mem[5431];

   memory[1358][0] = temp_mem[5432];
   memory[1358][1] = temp_mem[5433];
   memory[1358][2] = temp_mem[5434];
   memory[1358][3] = temp_mem[5435];

   memory[1359][0] = temp_mem[5436];
   memory[1359][1] = temp_mem[5437];
   memory[1359][2] = temp_mem[5438];
   memory[1359][3] = temp_mem[5439];

   memory[1360][0] = temp_mem[5440];
   memory[1360][1] = temp_mem[5441];
   memory[1360][2] = temp_mem[5442];
   memory[1360][3] = temp_mem[5443];

   memory[1361][0] = temp_mem[5444];
   memory[1361][1] = temp_mem[5445];
   memory[1361][2] = temp_mem[5446];
   memory[1361][3] = temp_mem[5447];

   memory[1362][0] = temp_mem[5448];
   memory[1362][1] = temp_mem[5449];
   memory[1362][2] = temp_mem[5450];
   memory[1362][3] = temp_mem[5451];

   memory[1363][0] = temp_mem[5452];
   memory[1363][1] = temp_mem[5453];
   memory[1363][2] = temp_mem[5454];
   memory[1363][3] = temp_mem[5455];

   memory[1364][0] = temp_mem[5456];
   memory[1364][1] = temp_mem[5457];
   memory[1364][2] = temp_mem[5458];
   memory[1364][3] = temp_mem[5459];

   memory[1365][0] = temp_mem[5460];
   memory[1365][1] = temp_mem[5461];
   memory[1365][2] = temp_mem[5462];
   memory[1365][3] = temp_mem[5463];

   memory[1366][0] = temp_mem[5464];
   memory[1366][1] = temp_mem[5465];
   memory[1366][2] = temp_mem[5466];
   memory[1366][3] = temp_mem[5467];

   memory[1367][0] = temp_mem[5468];
   memory[1367][1] = temp_mem[5469];
   memory[1367][2] = temp_mem[5470];
   memory[1367][3] = temp_mem[5471];

   memory[1368][0] = temp_mem[5472];
   memory[1368][1] = temp_mem[5473];
   memory[1368][2] = temp_mem[5474];
   memory[1368][3] = temp_mem[5475];

   memory[1369][0] = temp_mem[5476];
   memory[1369][1] = temp_mem[5477];
   memory[1369][2] = temp_mem[5478];
   memory[1369][3] = temp_mem[5479];

   memory[1370][0] = temp_mem[5480];
   memory[1370][1] = temp_mem[5481];
   memory[1370][2] = temp_mem[5482];
   memory[1370][3] = temp_mem[5483];

   memory[1371][0] = temp_mem[5484];
   memory[1371][1] = temp_mem[5485];
   memory[1371][2] = temp_mem[5486];
   memory[1371][3] = temp_mem[5487];

   memory[1372][0] = temp_mem[5488];
   memory[1372][1] = temp_mem[5489];
   memory[1372][2] = temp_mem[5490];
   memory[1372][3] = temp_mem[5491];

   memory[1373][0] = temp_mem[5492];
   memory[1373][1] = temp_mem[5493];
   memory[1373][2] = temp_mem[5494];
   memory[1373][3] = temp_mem[5495];

   memory[1374][0] = temp_mem[5496];
   memory[1374][1] = temp_mem[5497];
   memory[1374][2] = temp_mem[5498];
   memory[1374][3] = temp_mem[5499];

   memory[1375][0] = temp_mem[5500];
   memory[1375][1] = temp_mem[5501];
   memory[1375][2] = temp_mem[5502];
   memory[1375][3] = temp_mem[5503];

   memory[1376][0] = temp_mem[5504];
   memory[1376][1] = temp_mem[5505];
   memory[1376][2] = temp_mem[5506];
   memory[1376][3] = temp_mem[5507];

   memory[1377][0] = temp_mem[5508];
   memory[1377][1] = temp_mem[5509];
   memory[1377][2] = temp_mem[5510];
   memory[1377][3] = temp_mem[5511];

   memory[1378][0] = temp_mem[5512];
   memory[1378][1] = temp_mem[5513];
   memory[1378][2] = temp_mem[5514];
   memory[1378][3] = temp_mem[5515];

   memory[1379][0] = temp_mem[5516];
   memory[1379][1] = temp_mem[5517];
   memory[1379][2] = temp_mem[5518];
   memory[1379][3] = temp_mem[5519];

   memory[1380][0] = temp_mem[5520];
   memory[1380][1] = temp_mem[5521];
   memory[1380][2] = temp_mem[5522];
   memory[1380][3] = temp_mem[5523];

   memory[1381][0] = temp_mem[5524];
   memory[1381][1] = temp_mem[5525];
   memory[1381][2] = temp_mem[5526];
   memory[1381][3] = temp_mem[5527];

   memory[1382][0] = temp_mem[5528];
   memory[1382][1] = temp_mem[5529];
   memory[1382][2] = temp_mem[5530];
   memory[1382][3] = temp_mem[5531];

   memory[1383][0] = temp_mem[5532];
   memory[1383][1] = temp_mem[5533];
   memory[1383][2] = temp_mem[5534];
   memory[1383][3] = temp_mem[5535];

   memory[1384][0] = temp_mem[5536];
   memory[1384][1] = temp_mem[5537];
   memory[1384][2] = temp_mem[5538];
   memory[1384][3] = temp_mem[5539];

   memory[1385][0] = temp_mem[5540];
   memory[1385][1] = temp_mem[5541];
   memory[1385][2] = temp_mem[5542];
   memory[1385][3] = temp_mem[5543];

   memory[1386][0] = temp_mem[5544];
   memory[1386][1] = temp_mem[5545];
   memory[1386][2] = temp_mem[5546];
   memory[1386][3] = temp_mem[5547];

   memory[1387][0] = temp_mem[5548];
   memory[1387][1] = temp_mem[5549];
   memory[1387][2] = temp_mem[5550];
   memory[1387][3] = temp_mem[5551];

   memory[1388][0] = temp_mem[5552];
   memory[1388][1] = temp_mem[5553];
   memory[1388][2] = temp_mem[5554];
   memory[1388][3] = temp_mem[5555];

   memory[1389][0] = temp_mem[5556];
   memory[1389][1] = temp_mem[5557];
   memory[1389][2] = temp_mem[5558];
   memory[1389][3] = temp_mem[5559];

   memory[1390][0] = temp_mem[5560];
   memory[1390][1] = temp_mem[5561];
   memory[1390][2] = temp_mem[5562];
   memory[1390][3] = temp_mem[5563];

   memory[1391][0] = temp_mem[5564];
   memory[1391][1] = temp_mem[5565];
   memory[1391][2] = temp_mem[5566];
   memory[1391][3] = temp_mem[5567];

   memory[1392][0] = temp_mem[5568];
   memory[1392][1] = temp_mem[5569];
   memory[1392][2] = temp_mem[5570];
   memory[1392][3] = temp_mem[5571];

   memory[1393][0] = temp_mem[5572];
   memory[1393][1] = temp_mem[5573];
   memory[1393][2] = temp_mem[5574];
   memory[1393][3] = temp_mem[5575];

   memory[1394][0] = temp_mem[5576];
   memory[1394][1] = temp_mem[5577];
   memory[1394][2] = temp_mem[5578];
   memory[1394][3] = temp_mem[5579];

   memory[1395][0] = temp_mem[5580];
   memory[1395][1] = temp_mem[5581];
   memory[1395][2] = temp_mem[5582];
   memory[1395][3] = temp_mem[5583];

   memory[1396][0] = temp_mem[5584];
   memory[1396][1] = temp_mem[5585];
   memory[1396][2] = temp_mem[5586];
   memory[1396][3] = temp_mem[5587];

   memory[1397][0] = temp_mem[5588];
   memory[1397][1] = temp_mem[5589];
   memory[1397][2] = temp_mem[5590];
   memory[1397][3] = temp_mem[5591];

   memory[1398][0] = temp_mem[5592];
   memory[1398][1] = temp_mem[5593];
   memory[1398][2] = temp_mem[5594];
   memory[1398][3] = temp_mem[5595];

   memory[1399][0] = temp_mem[5596];
   memory[1399][1] = temp_mem[5597];
   memory[1399][2] = temp_mem[5598];
   memory[1399][3] = temp_mem[5599];

   memory[1400][0] = temp_mem[5600];
   memory[1400][1] = temp_mem[5601];
   memory[1400][2] = temp_mem[5602];
   memory[1400][3] = temp_mem[5603];

   memory[1401][0] = temp_mem[5604];
   memory[1401][1] = temp_mem[5605];
   memory[1401][2] = temp_mem[5606];
   memory[1401][3] = temp_mem[5607];

   memory[1402][0] = temp_mem[5608];
   memory[1402][1] = temp_mem[5609];
   memory[1402][2] = temp_mem[5610];
   memory[1402][3] = temp_mem[5611];

   memory[1403][0] = temp_mem[5612];
   memory[1403][1] = temp_mem[5613];
   memory[1403][2] = temp_mem[5614];
   memory[1403][3] = temp_mem[5615];

   memory[1404][0] = temp_mem[5616];
   memory[1404][1] = temp_mem[5617];
   memory[1404][2] = temp_mem[5618];
   memory[1404][3] = temp_mem[5619];

   memory[1405][0] = temp_mem[5620];
   memory[1405][1] = temp_mem[5621];
   memory[1405][2] = temp_mem[5622];
   memory[1405][3] = temp_mem[5623];

   memory[1406][0] = temp_mem[5624];
   memory[1406][1] = temp_mem[5625];
   memory[1406][2] = temp_mem[5626];
   memory[1406][3] = temp_mem[5627];

   memory[1407][0] = temp_mem[5628];
   memory[1407][1] = temp_mem[5629];
   memory[1407][2] = temp_mem[5630];
   memory[1407][3] = temp_mem[5631];

   memory[1408][0] = temp_mem[5632];
   memory[1408][1] = temp_mem[5633];
   memory[1408][2] = temp_mem[5634];
   memory[1408][3] = temp_mem[5635];

   memory[1409][0] = temp_mem[5636];
   memory[1409][1] = temp_mem[5637];
   memory[1409][2] = temp_mem[5638];
   memory[1409][3] = temp_mem[5639];

   memory[1410][0] = temp_mem[5640];
   memory[1410][1] = temp_mem[5641];
   memory[1410][2] = temp_mem[5642];
   memory[1410][3] = temp_mem[5643];

   memory[1411][0] = temp_mem[5644];
   memory[1411][1] = temp_mem[5645];
   memory[1411][2] = temp_mem[5646];
   memory[1411][3] = temp_mem[5647];

   memory[1412][0] = temp_mem[5648];
   memory[1412][1] = temp_mem[5649];
   memory[1412][2] = temp_mem[5650];
   memory[1412][3] = temp_mem[5651];

   memory[1413][0] = temp_mem[5652];
   memory[1413][1] = temp_mem[5653];
   memory[1413][2] = temp_mem[5654];
   memory[1413][3] = temp_mem[5655];

   memory[1414][0] = temp_mem[5656];
   memory[1414][1] = temp_mem[5657];
   memory[1414][2] = temp_mem[5658];
   memory[1414][3] = temp_mem[5659];

   memory[1415][0] = temp_mem[5660];
   memory[1415][1] = temp_mem[5661];
   memory[1415][2] = temp_mem[5662];
   memory[1415][3] = temp_mem[5663];

   memory[1416][0] = temp_mem[5664];
   memory[1416][1] = temp_mem[5665];
   memory[1416][2] = temp_mem[5666];
   memory[1416][3] = temp_mem[5667];

   memory[1417][0] = temp_mem[5668];
   memory[1417][1] = temp_mem[5669];
   memory[1417][2] = temp_mem[5670];
   memory[1417][3] = temp_mem[5671];

   memory[1418][0] = temp_mem[5672];
   memory[1418][1] = temp_mem[5673];
   memory[1418][2] = temp_mem[5674];
   memory[1418][3] = temp_mem[5675];

   memory[1419][0] = temp_mem[5676];
   memory[1419][1] = temp_mem[5677];
   memory[1419][2] = temp_mem[5678];
   memory[1419][3] = temp_mem[5679];

   memory[1420][0] = temp_mem[5680];
   memory[1420][1] = temp_mem[5681];
   memory[1420][2] = temp_mem[5682];
   memory[1420][3] = temp_mem[5683];

   memory[1421][0] = temp_mem[5684];
   memory[1421][1] = temp_mem[5685];
   memory[1421][2] = temp_mem[5686];
   memory[1421][3] = temp_mem[5687];

   memory[1422][0] = temp_mem[5688];
   memory[1422][1] = temp_mem[5689];
   memory[1422][2] = temp_mem[5690];
   memory[1422][3] = temp_mem[5691];

   memory[1423][0] = temp_mem[5692];
   memory[1423][1] = temp_mem[5693];
   memory[1423][2] = temp_mem[5694];
   memory[1423][3] = temp_mem[5695];

   memory[1424][0] = temp_mem[5696];
   memory[1424][1] = temp_mem[5697];
   memory[1424][2] = temp_mem[5698];
   memory[1424][3] = temp_mem[5699];

   memory[1425][0] = temp_mem[5700];
   memory[1425][1] = temp_mem[5701];
   memory[1425][2] = temp_mem[5702];
   memory[1425][3] = temp_mem[5703];

   memory[1426][0] = temp_mem[5704];
   memory[1426][1] = temp_mem[5705];
   memory[1426][2] = temp_mem[5706];
   memory[1426][3] = temp_mem[5707];

   memory[1427][0] = temp_mem[5708];
   memory[1427][1] = temp_mem[5709];
   memory[1427][2] = temp_mem[5710];
   memory[1427][3] = temp_mem[5711];

   memory[1428][0] = temp_mem[5712];
   memory[1428][1] = temp_mem[5713];
   memory[1428][2] = temp_mem[5714];
   memory[1428][3] = temp_mem[5715];

   memory[1429][0] = temp_mem[5716];
   memory[1429][1] = temp_mem[5717];
   memory[1429][2] = temp_mem[5718];
   memory[1429][3] = temp_mem[5719];

   memory[1430][0] = temp_mem[5720];
   memory[1430][1] = temp_mem[5721];
   memory[1430][2] = temp_mem[5722];
   memory[1430][3] = temp_mem[5723];

   memory[1431][0] = temp_mem[5724];
   memory[1431][1] = temp_mem[5725];
   memory[1431][2] = temp_mem[5726];
   memory[1431][3] = temp_mem[5727];

   memory[1432][0] = temp_mem[5728];
   memory[1432][1] = temp_mem[5729];
   memory[1432][2] = temp_mem[5730];
   memory[1432][3] = temp_mem[5731];

   memory[1433][0] = temp_mem[5732];
   memory[1433][1] = temp_mem[5733];
   memory[1433][2] = temp_mem[5734];
   memory[1433][3] = temp_mem[5735];

   memory[1434][0] = temp_mem[5736];
   memory[1434][1] = temp_mem[5737];
   memory[1434][2] = temp_mem[5738];
   memory[1434][3] = temp_mem[5739];

   memory[1435][0] = temp_mem[5740];
   memory[1435][1] = temp_mem[5741];
   memory[1435][2] = temp_mem[5742];
   memory[1435][3] = temp_mem[5743];

   memory[1436][0] = temp_mem[5744];
   memory[1436][1] = temp_mem[5745];
   memory[1436][2] = temp_mem[5746];
   memory[1436][3] = temp_mem[5747];

   memory[1437][0] = temp_mem[5748];
   memory[1437][1] = temp_mem[5749];
   memory[1437][2] = temp_mem[5750];
   memory[1437][3] = temp_mem[5751];

   memory[1438][0] = temp_mem[5752];
   memory[1438][1] = temp_mem[5753];
   memory[1438][2] = temp_mem[5754];
   memory[1438][3] = temp_mem[5755];

   memory[1439][0] = temp_mem[5756];
   memory[1439][1] = temp_mem[5757];
   memory[1439][2] = temp_mem[5758];
   memory[1439][3] = temp_mem[5759];

   memory[1440][0] = temp_mem[5760];
   memory[1440][1] = temp_mem[5761];
   memory[1440][2] = temp_mem[5762];
   memory[1440][3] = temp_mem[5763];

   memory[1441][0] = temp_mem[5764];
   memory[1441][1] = temp_mem[5765];
   memory[1441][2] = temp_mem[5766];
   memory[1441][3] = temp_mem[5767];

   memory[1442][0] = temp_mem[5768];
   memory[1442][1] = temp_mem[5769];
   memory[1442][2] = temp_mem[5770];
   memory[1442][3] = temp_mem[5771];

   memory[1443][0] = temp_mem[5772];
   memory[1443][1] = temp_mem[5773];
   memory[1443][2] = temp_mem[5774];
   memory[1443][3] = temp_mem[5775];

   memory[1444][0] = temp_mem[5776];
   memory[1444][1] = temp_mem[5777];
   memory[1444][2] = temp_mem[5778];
   memory[1444][3] = temp_mem[5779];

   memory[1445][0] = temp_mem[5780];
   memory[1445][1] = temp_mem[5781];
   memory[1445][2] = temp_mem[5782];
   memory[1445][3] = temp_mem[5783];

   memory[1446][0] = temp_mem[5784];
   memory[1446][1] = temp_mem[5785];
   memory[1446][2] = temp_mem[5786];
   memory[1446][3] = temp_mem[5787];

   memory[1447][0] = temp_mem[5788];
   memory[1447][1] = temp_mem[5789];
   memory[1447][2] = temp_mem[5790];
   memory[1447][3] = temp_mem[5791];

   memory[1448][0] = temp_mem[5792];
   memory[1448][1] = temp_mem[5793];
   memory[1448][2] = temp_mem[5794];
   memory[1448][3] = temp_mem[5795];

   memory[1449][0] = temp_mem[5796];
   memory[1449][1] = temp_mem[5797];
   memory[1449][2] = temp_mem[5798];
   memory[1449][3] = temp_mem[5799];
	
	memory[1450][0] = temp_mem[5800];
   memory[1450][1] = temp_mem[5801];
   memory[1450][2] = temp_mem[5802];
   memory[1450][3] = temp_mem[5803];

	memory[1451][0] = temp_mem[5804];
	memory[1451][1] = temp_mem[5805];
	memory[1451][2] = temp_mem[5806];
	memory[1451][3] = temp_mem[5807];

	memory[1452][0] = temp_mem[5808];
	memory[1452][1] = temp_mem[5809];
	memory[1452][2] = temp_mem[5810];
	memory[1452][3] = temp_mem[5811];

	memory[1453][0] = temp_mem[5812];
	memory[1453][1] = temp_mem[5813];
	memory[1453][2] = temp_mem[5814];
	memory[1453][3] = temp_mem[5815];

	memory[1454][0] = temp_mem[5816];
	memory[1454][1] = temp_mem[5817];
	memory[1454][2] = temp_mem[5818];
	memory[1454][3] = temp_mem[5819];

	memory[1455][0] = temp_mem[5820];
	memory[1455][1] = temp_mem[5821];
	memory[1455][2] = temp_mem[5822];
	memory[1455][3] = temp_mem[5823];

	memory[1456][0] = temp_mem[5824];
	memory[1456][1] = temp_mem[5825];
	memory[1456][2] = temp_mem[5826];
	memory[1456][3] = temp_mem[5827];

	memory[1457][0] = temp_mem[5828];
	memory[1457][1] = temp_mem[5829];
	memory[1457][2] = temp_mem[5830];
	memory[1457][3] = temp_mem[5831];

	memory[1458][0] = temp_mem[5832];
	memory[1458][1] = temp_mem[5833];
	memory[1458][2] = temp_mem[5834];
	memory[1458][3] = temp_mem[5835];

	memory[1459][0] = temp_mem[5836];
	memory[1459][1] = temp_mem[5837];
	memory[1459][2] = temp_mem[5838];
	memory[1459][3] = temp_mem[5839];

	memory[1460][0] = temp_mem[5840];
	memory[1460][1] = temp_mem[5841];
	memory[1460][2] = temp_mem[5842];
	memory[1460][3] = temp_mem[5843];

	memory[1461][0] = temp_mem[5844];
	memory[1461][1] = temp_mem[5845];
	memory[1461][2] = temp_mem[5846];
	memory[1461][3] = temp_mem[5847];

	memory[1462][0] = temp_mem[5848];
	memory[1462][1] = temp_mem[5849];
	memory[1462][2] = temp_mem[5850];
	memory[1462][3] = temp_mem[5851];

	memory[1463][0] = temp_mem[5852];
	memory[1463][1] = temp_mem[5853];
	memory[1463][2] = temp_mem[5854];
	memory[1463][3] = temp_mem[5855];

	memory[1464][0] = temp_mem[5856];
	memory[1464][1] = temp_mem[5857];
	memory[1464][2] = temp_mem[5858];
	memory[1464][3] = temp_mem[5859];

	memory[1465][0] = temp_mem[5860];
	memory[1465][1] = temp_mem[5861];
	memory[1465][2] = temp_mem[5862];
	memory[1465][3] = temp_mem[5863];

	memory[1466][0] = temp_mem[5864];
	memory[1466][1] = temp_mem[5865];
	memory[1466][2] = temp_mem[5866];
	memory[1466][3] = temp_mem[5867];

	memory[1467][0] = temp_mem[5868];
	memory[1467][1] = temp_mem[5869];
	memory[1467][2] = temp_mem[5870];
	memory[1467][3] = temp_mem[5871];

	memory[1468][0] = temp_mem[5872];
	memory[1468][1] = temp_mem[5873];
	memory[1468][2] = temp_mem[5874];
	memory[1468][3] = temp_mem[5875];

	memory[1469][0] = temp_mem[5876];
	memory[1469][1] = temp_mem[5877];
	memory[1469][2] = temp_mem[5878];
	memory[1469][3] = temp_mem[5879];

	memory[1470][0] = temp_mem[5880];
	memory[1470][1] = temp_mem[5881];
	memory[1470][2] = temp_mem[5882];
	memory[1470][3] = temp_mem[5883];

	memory[1471][0] = temp_mem[5884];
	memory[1471][1] = temp_mem[5885];
	memory[1471][2] = temp_mem[5886];
	memory[1471][3] = temp_mem[5887];

	memory[1472][0] = temp_mem[5888];
	memory[1472][1] = temp_mem[5889];
	memory[1472][2] = temp_mem[5890];
	memory[1472][3] = temp_mem[5891];

	memory[1473][0] = temp_mem[5892];
	memory[1473][1] = temp_mem[5893];
	memory[1473][2] = temp_mem[5894];
	memory[1473][3] = temp_mem[5895];

	memory[1474][0] = temp_mem[5896];
	memory[1474][1] = temp_mem[5897];
	memory[1474][2] = temp_mem[5898];
	memory[1474][3] = temp_mem[5899];

	memory[1475][0] = temp_mem[5900];
	memory[1475][1] = temp_mem[5901];
	memory[1475][2] = temp_mem[5902];
	memory[1475][3] = temp_mem[5903];

	memory[1476][0] = temp_mem[5904];
	memory[1476][1] = temp_mem[5905];
	memory[1476][2] = temp_mem[5906];
	memory[1476][3] = temp_mem[5907];

	memory[1477][0] = temp_mem[5908];
	memory[1477][1] = temp_mem[5909];
	memory[1477][2] = temp_mem[5910];
	memory[1477][3] = temp_mem[5911];

	memory[1478][0] = temp_mem[5912];
	memory[1478][1] = temp_mem[5913];
	memory[1478][2] = temp_mem[5914];
	memory[1478][3] = temp_mem[5915];

	memory[1479][0] = temp_mem[5916];
	memory[1479][1] = temp_mem[5917];
	memory[1479][2] = temp_mem[5918];
	memory[1479][3] = temp_mem[5919];

	memory[1480][0] = temp_mem[5920];
	memory[1480][1] = temp_mem[5921];
	memory[1480][2] = temp_mem[5922];
	memory[1480][3] = temp_mem[5923];

	memory[1481][0] = temp_mem[5924];
	memory[1481][1] = temp_mem[5925];
	memory[1481][2] = temp_mem[5926];
	memory[1481][3] = temp_mem[5927];

	memory[1482][0] = temp_mem[5928];
	memory[1482][1] = temp_mem[5929];
	memory[1482][2] = temp_mem[5930];
	memory[1482][3] = temp_mem[5931];

	memory[1483][0] = temp_mem[5932];
	memory[1483][1] = temp_mem[5933];
	memory[1483][2] = temp_mem[5934];
	memory[1483][3] = temp_mem[5935];

	memory[1484][0] = temp_mem[5936];
	memory[1484][1] = temp_mem[5937];
	memory[1484][2] = temp_mem[5938];
	memory[1484][3] = temp_mem[5939];

	memory[1485][0] = temp_mem[5940];
	memory[1485][1] = temp_mem[5941];
	memory[1485][2] = temp_mem[5942];
	memory[1485][3] = temp_mem[5943];

	memory[1486][0] = temp_mem[5944];
	memory[1486][1] = temp_mem[5945];
	memory[1486][2] = temp_mem[5946];
	memory[1486][3] = temp_mem[5947];

	memory[1487][0] = temp_mem[5948];
	memory[1487][1] = temp_mem[5949];
	memory[1487][2] = temp_mem[5950];
	memory[1487][3] = temp_mem[5951];

	memory[1488][0] = temp_mem[5952];
	memory[1488][1] = temp_mem[5953];
	memory[1488][2] = temp_mem[5954];
	memory[1488][3] = temp_mem[5955];

	memory[1489][0] = temp_mem[5956];
	memory[1489][1] = temp_mem[5957];
	memory[1489][2] = temp_mem[5958];
	memory[1489][3] = temp_mem[5959];

	memory[1490][0] = temp_mem[5960];
	memory[1490][1] = temp_mem[5961];
	memory[1490][2] = temp_mem[5962];
	memory[1490][3] = temp_mem[5963];

	memory[1491][0] = temp_mem[5964];
	memory[1491][1] = temp_mem[5965];
	memory[1491][2] = temp_mem[5966];
	memory[1491][3] = temp_mem[5967];

	memory[1492][0] = temp_mem[5968];
	memory[1492][1] = temp_mem[5969];
	memory[1492][2] = temp_mem[5970];
	memory[1492][3] = temp_mem[5971];

	memory[1493][0] = temp_mem[5972];
	memory[1493][1] = temp_mem[5973];
	memory[1493][2] = temp_mem[5974];
	memory[1493][3] = temp_mem[5975];

	memory[1494][0] = temp_mem[5976];
	memory[1494][1] = temp_mem[5977];
	memory[1494][2] = temp_mem[5978];
	memory[1494][3] = temp_mem[5979];

	memory[1495][0] = temp_mem[5980];
	memory[1495][1] = temp_mem[5981];
	memory[1495][2] = temp_mem[5982];
	memory[1495][3] = temp_mem[5983];

	memory[1496][0] = temp_mem[5984];
	memory[1496][1] = temp_mem[5985];
	memory[1496][2] = temp_mem[5986];
	memory[1496][3] = temp_mem[5987];

	memory[1497][0] = temp_mem[5988];
	memory[1497][1] = temp_mem[5989];
	memory[1497][2] = temp_mem[5990];
	memory[1497][3] = temp_mem[5991];

	memory[1498][0] = temp_mem[5992];
	memory[1498][1] = temp_mem[5993];
	memory[1498][2] = temp_mem[5994];
	memory[1498][3] = temp_mem[5995];

	memory[1499][0] = temp_mem[5996];
	memory[1499][1] = temp_mem[5997];
	memory[1499][2] = temp_mem[5998];
	memory[1499][3] = temp_mem[5999];

	memory[1500][0] = temp_mem[6000];
	memory[1500][1] = temp_mem[6001];
	memory[1500][2] = temp_mem[6002];
	memory[1500][3] = temp_mem[6003];

	memory[1501][0] = temp_mem[6004];
	memory[1501][1] = temp_mem[6005];
	memory[1501][2] = temp_mem[6006];
	memory[1501][3] = temp_mem[6007];

	memory[1502][0] = temp_mem[6008];
	memory[1502][1] = temp_mem[6009];
	memory[1502][2] = temp_mem[6010];
	memory[1502][3] = temp_mem[6011];

	memory[1503][0] = temp_mem[6012];
	memory[1503][1] = temp_mem[6013];
	memory[1503][2] = temp_mem[6014];
	memory[1503][3] = temp_mem[6015];

	memory[1504][0] = temp_mem[6016];
	memory[1504][1] = temp_mem[6017];
	memory[1504][2] = temp_mem[6018];
	memory[1504][3] = temp_mem[6019];

	memory[1505][0] = temp_mem[6020];
	memory[1505][1] = temp_mem[6021];
	memory[1505][2] = temp_mem[6022];
	memory[1505][3] = temp_mem[6023];

	memory[1506][0] = temp_mem[6024];
	memory[1506][1] = temp_mem[6025];
	memory[1506][2] = temp_mem[6026];
	memory[1506][3] = temp_mem[6027];

	memory[1507][0] = temp_mem[6028];
	memory[1507][1] = temp_mem[6029];
	memory[1507][2] = temp_mem[6030];
	memory[1507][3] = temp_mem[6031];

	memory[1508][0] = temp_mem[6032];
	memory[1508][1] = temp_mem[6033];
	memory[1508][2] = temp_mem[6034];
	memory[1508][3] = temp_mem[6035];

	memory[1509][0] = temp_mem[6036];
	memory[1509][1] = temp_mem[6037];
	memory[1509][2] = temp_mem[6038];
	memory[1509][3] = temp_mem[6039];

	memory[1510][0] = temp_mem[6040];
	memory[1510][1] = temp_mem[6041];
	memory[1510][2] = temp_mem[6042];
	memory[1510][3] = temp_mem[6043];

	memory[1511][0] = temp_mem[6044];
	memory[1511][1] = temp_mem[6045];
	memory[1511][2] = temp_mem[6046];
	memory[1511][3] = temp_mem[6047];

	memory[1512][0] = temp_mem[6048];
	memory[1512][1] = temp_mem[6049];
	memory[1512][2] = temp_mem[6050];
	memory[1512][3] = temp_mem[6051];

	memory[1513][0] = temp_mem[6052];
	memory[1513][1] = temp_mem[6053];
	memory[1513][2] = temp_mem[6054];
	memory[1513][3] = temp_mem[6055];

	memory[1514][0] = temp_mem[6056];
	memory[1514][1] = temp_mem[6057];
	memory[1514][2] = temp_mem[6058];
	memory[1514][3] = temp_mem[6059];

	memory[1515][0] = temp_mem[6060];
	memory[1515][1] = temp_mem[6061];
	memory[1515][2] = temp_mem[6062];
	memory[1515][3] = temp_mem[6063];

	memory[1516][0] = temp_mem[6064];
	memory[1516][1] = temp_mem[6065];
	memory[1516][2] = temp_mem[6066];
	memory[1516][3] = temp_mem[6067];

	memory[1517][0] = temp_mem[6068];
	memory[1517][1] = temp_mem[6069];
	memory[1517][2] = temp_mem[6070];
	memory[1517][3] = temp_mem[6071];

	memory[1518][0] = temp_mem[6072];
	memory[1518][1] = temp_mem[6073];
	memory[1518][2] = temp_mem[6074];
	memory[1518][3] = temp_mem[6075];

	memory[1519][0] = temp_mem[6076];
	memory[1519][1] = temp_mem[6077];
	memory[1519][2] = temp_mem[6078];
	memory[1519][3] = temp_mem[6079];

	memory[1520][0] = temp_mem[6080];
	memory[1520][1] = temp_mem[6081];
	memory[1520][2] = temp_mem[6082];
	memory[1520][3] = temp_mem[6083];

	memory[1521][0] = temp_mem[6084];
	memory[1521][1] = temp_mem[6085];
	memory[1521][2] = temp_mem[6086];
	memory[1521][3] = temp_mem[6087];

	memory[1522][0] = temp_mem[6088];
	memory[1522][1] = temp_mem[6089];
	memory[1522][2] = temp_mem[6090];
	memory[1522][3] = temp_mem[6091];

	memory[1523][0] = temp_mem[6092];
	memory[1523][1] = temp_mem[6093];
	memory[1523][2] = temp_mem[6094];
	memory[1523][3] = temp_mem[6095];

	memory[1524][0] = temp_mem[6096];
	memory[1524][1] = temp_mem[6097];
	memory[1524][2] = temp_mem[6098];
	memory[1524][3] = temp_mem[6099];

	memory[1525][0] = temp_mem[6100];
	memory[1525][1] = temp_mem[6101];
	memory[1525][2] = temp_mem[6102];
	memory[1525][3] = temp_mem[6103];

	memory[1526][0] = temp_mem[6104];
	memory[1526][1] = temp_mem[6105];
	memory[1526][2] = temp_mem[6106];
	memory[1526][3] = temp_mem[6107];

	memory[1527][0] = temp_mem[6108];
	memory[1527][1] = temp_mem[6109];
	memory[1527][2] = temp_mem[6110];
	memory[1527][3] = temp_mem[6111];

	memory[1528][0] = temp_mem[6112];
	memory[1528][1] = temp_mem[6113];
	memory[1528][2] = temp_mem[6114];
	memory[1528][3] = temp_mem[6115];

	memory[1529][0] = temp_mem[6116];
	memory[1529][1] = temp_mem[6117];
	memory[1529][2] = temp_mem[6118];
	memory[1529][3] = temp_mem[6119];

	memory[1530][0] = temp_mem[6120];
	memory[1530][1] = temp_mem[6121];
	memory[1530][2] = temp_mem[6122];
	memory[1530][3] = temp_mem[6123];

	memory[1531][0] = temp_mem[6124];
	memory[1531][1] = temp_mem[6125];
	memory[1531][2] = temp_mem[6126];
	memory[1531][3] = temp_mem[6127];

	memory[1532][0] = temp_mem[6128];
	memory[1532][1] = temp_mem[6129];
	memory[1532][2] = temp_mem[6130];
	memory[1532][3] = temp_mem[6131];

	memory[1533][0] = temp_mem[6132];
	memory[1533][1] = temp_mem[6133];
	memory[1533][2] = temp_mem[6134];
	memory[1533][3] = temp_mem[6135];

	memory[1534][0] = temp_mem[6136];
	memory[1534][1] = temp_mem[6137];
	memory[1534][2] = temp_mem[6138];
	memory[1534][3] = temp_mem[6139];

	memory[1535][0] = temp_mem[6140];
	memory[1535][1] = temp_mem[6141];
	memory[1535][2] = temp_mem[6142];
	memory[1535][3] = temp_mem[6143];

	memory[1536][0] = temp_mem[6144];
	memory[1536][1] = temp_mem[6145];
	memory[1536][2] = temp_mem[6146];
	memory[1536][3] = temp_mem[6147];

	memory[1537][0] = temp_mem[6148];
	memory[1537][1] = temp_mem[6149];
	memory[1537][2] = temp_mem[6150];
	memory[1537][3] = temp_mem[6151];

	memory[1538][0] = temp_mem[6152];
	memory[1538][1] = temp_mem[6153];
	memory[1538][2] = temp_mem[6154];
	memory[1538][3] = temp_mem[6155];

	memory[1539][0] = temp_mem[6156];
	memory[1539][1] = temp_mem[6157];
	memory[1539][2] = temp_mem[6158];
	memory[1539][3] = temp_mem[6159];

	memory[1540][0] = temp_mem[6160];
	memory[1540][1] = temp_mem[6161];
	memory[1540][2] = temp_mem[6162];
	memory[1540][3] = temp_mem[6163];

	memory[1541][0] = temp_mem[6164];
	memory[1541][1] = temp_mem[6165];
	memory[1541][2] = temp_mem[6166];
	memory[1541][3] = temp_mem[6167];

	memory[1542][0] = temp_mem[6168];
	memory[1542][1] = temp_mem[6169];
	memory[1542][2] = temp_mem[6170];
	memory[1542][3] = temp_mem[6171];

	memory[1543][0] = temp_mem[6172];
	memory[1543][1] = temp_mem[6173];
	memory[1543][2] = temp_mem[6174];
	memory[1543][3] = temp_mem[6175];

	memory[1544][0] = temp_mem[6176];
	memory[1544][1] = temp_mem[6177];
	memory[1544][2] = temp_mem[6178];
	memory[1544][3] = temp_mem[6179];

	memory[1545][0] = temp_mem[6180];
	memory[1545][1] = temp_mem[6181];
	memory[1545][2] = temp_mem[6182];
	memory[1545][3] = temp_mem[6183];

	memory[1546][0] = temp_mem[6184];
	memory[1546][1] = temp_mem[6185];
	memory[1546][2] = temp_mem[6186];
	memory[1546][3] = temp_mem[6187];

	memory[1547][0] = temp_mem[6188];
	memory[1547][1] = temp_mem[6189];
	memory[1547][2] = temp_mem[6190];
	memory[1547][3] = temp_mem[6191];

	memory[1548][0] = temp_mem[6192];
	memory[1548][1] = temp_mem[6193];
	memory[1548][2] = temp_mem[6194];
	memory[1548][3] = temp_mem[6195];

	memory[1549][0] = temp_mem[6196];
	memory[1549][1] = temp_mem[6197];
	memory[1549][2] = temp_mem[6198];
	memory[1549][3] = temp_mem[6199];

	memory[1550][0] = temp_mem[6200];
	memory[1550][1] = temp_mem[6201];
	memory[1550][2] = temp_mem[6202];
	memory[1550][3] = temp_mem[6203];

	memory[1551][0] = temp_mem[6204];
	memory[1551][1] = temp_mem[6205];
	memory[1551][2] = temp_mem[6206];
	memory[1551][3] = temp_mem[6207];

	memory[1552][0] = temp_mem[6208];
	memory[1552][1] = temp_mem[6209];
	memory[1552][2] = temp_mem[6210];
	memory[1552][3] = temp_mem[6211];

	memory[1553][0] = temp_mem[6212];
	memory[1553][1] = temp_mem[6213];
	memory[1553][2] = temp_mem[6214];
	memory[1553][3] = temp_mem[6215];

	memory[1554][0] = temp_mem[6216];
	memory[1554][1] = temp_mem[6217];
	memory[1554][2] = temp_mem[6218];
	memory[1554][3] = temp_mem[6219];

	memory[1555][0] = temp_mem[6220];
	memory[1555][1] = temp_mem[6221];
	memory[1555][2] = temp_mem[6222];
	memory[1555][3] = temp_mem[6223];

	memory[1556][0] = temp_mem[6224];
	memory[1556][1] = temp_mem[6225];
	memory[1556][2] = temp_mem[6226];
	memory[1556][3] = temp_mem[6227];

	memory[1557][0] = temp_mem[6228];
	memory[1557][1] = temp_mem[6229];
	memory[1557][2] = temp_mem[6230];
	memory[1557][3] = temp_mem[6231];

	memory[1558][0] = temp_mem[6232];
	memory[1558][1] = temp_mem[6233];
	memory[1558][2] = temp_mem[6234];
	memory[1558][3] = temp_mem[6235];

	memory[1559][0] = temp_mem[6236];
	memory[1559][1] = temp_mem[6237];
	memory[1559][2] = temp_mem[6238];
	memory[1559][3] = temp_mem[6239];

	memory[1560][0] = temp_mem[6240];
	memory[1560][1] = temp_mem[6241];
	memory[1560][2] = temp_mem[6242];
	memory[1560][3] = temp_mem[6243];

	memory[1561][0] = temp_mem[6244];
	memory[1561][1] = temp_mem[6245];
	memory[1561][2] = temp_mem[6246];
	memory[1561][3] = temp_mem[6247];

	memory[1562][0] = temp_mem[6248];
	memory[1562][1] = temp_mem[6249];
	memory[1562][2] = temp_mem[6250];
	memory[1562][3] = temp_mem[6251];

	memory[1563][0] = temp_mem[6252];
	memory[1563][1] = temp_mem[6253];
	memory[1563][2] = temp_mem[6254];
	memory[1563][3] = temp_mem[6255];

	memory[1564][0] = temp_mem[6256];
	memory[1564][1] = temp_mem[6257];
	memory[1564][2] = temp_mem[6258];
	memory[1564][3] = temp_mem[6259];

	memory[1565][0] = temp_mem[6260];
	memory[1565][1] = temp_mem[6261];
	memory[1565][2] = temp_mem[6262];
	memory[1565][3] = temp_mem[6263];

	memory[1566][0] = temp_mem[6264];
	memory[1566][1] = temp_mem[6265];
	memory[1566][2] = temp_mem[6266];
	memory[1566][3] = temp_mem[6267];

	memory[1567][0] = temp_mem[6268];
	memory[1567][1] = temp_mem[6269];
	memory[1567][2] = temp_mem[6270];
	memory[1567][3] = temp_mem[6271];

	memory[1568][0] = temp_mem[6272];
	memory[1568][1] = temp_mem[6273];
	memory[1568][2] = temp_mem[6274];
	memory[1568][3] = temp_mem[6275];

	memory[1569][0] = temp_mem[6276];
	memory[1569][1] = temp_mem[6277];
	memory[1569][2] = temp_mem[6278];
	memory[1569][3] = temp_mem[6279];

	memory[1570][0] = temp_mem[6280];
	memory[1570][1] = temp_mem[6281];
	memory[1570][2] = temp_mem[6282];
	memory[1570][3] = temp_mem[6283];

	memory[1571][0] = temp_mem[6284];
	memory[1571][1] = temp_mem[6285];
	memory[1571][2] = temp_mem[6286];
	memory[1571][3] = temp_mem[6287];

	memory[1572][0] = temp_mem[6288];
	memory[1572][1] = temp_mem[6289];
	memory[1572][2] = temp_mem[6290];
	memory[1572][3] = temp_mem[6291];

	memory[1573][0] = temp_mem[6292];
	memory[1573][1] = temp_mem[6293];
	memory[1573][2] = temp_mem[6294];
	memory[1573][3] = temp_mem[6295];

	memory[1574][0] = temp_mem[6296];
	memory[1574][1] = temp_mem[6297];
	memory[1574][2] = temp_mem[6298];
	memory[1574][3] = temp_mem[6299];

	memory[1575][0] = temp_mem[6300];
	memory[1575][1] = temp_mem[6301];
	memory[1575][2] = temp_mem[6302];
	memory[1575][3] = temp_mem[6303];

	memory[1576][0] = temp_mem[6304];
	memory[1576][1] = temp_mem[6305];
	memory[1576][2] = temp_mem[6306];
	memory[1576][3] = temp_mem[6307];

	memory[1577][0] = temp_mem[6308];
	memory[1577][1] = temp_mem[6309];
	memory[1577][2] = temp_mem[6310];
	memory[1577][3] = temp_mem[6311];

	memory[1578][0] = temp_mem[6312];
	memory[1578][1] = temp_mem[6313];
	memory[1578][2] = temp_mem[6314];
	memory[1578][3] = temp_mem[6315];

	memory[1579][0] = temp_mem[6316];
	memory[1579][1] = temp_mem[6317];
	memory[1579][2] = temp_mem[6318];
	memory[1579][3] = temp_mem[6319];

	memory[1580][0] = temp_mem[6320];
	memory[1580][1] = temp_mem[6321];
	memory[1580][2] = temp_mem[6322];
	memory[1580][3] = temp_mem[6323];

	memory[1581][0] = temp_mem[6324];
	memory[1581][1] = temp_mem[6325];
	memory[1581][2] = temp_mem[6326];
	memory[1581][3] = temp_mem[6327];

	memory[1582][0] = temp_mem[6328];
	memory[1582][1] = temp_mem[6329];
	memory[1582][2] = temp_mem[6330];
	memory[1582][3] = temp_mem[6331];

	memory[1583][0] = temp_mem[6332];
	memory[1583][1] = temp_mem[6333];
	memory[1583][2] = temp_mem[6334];
	memory[1583][3] = temp_mem[6335];

	memory[1584][0] = temp_mem[6336];
	memory[1584][1] = temp_mem[6337];
	memory[1584][2] = temp_mem[6338];
	memory[1584][3] = temp_mem[6339];

	memory[1585][0] = temp_mem[6340];
	memory[1585][1] = temp_mem[6341];
	memory[1585][2] = temp_mem[6342];
	memory[1585][3] = temp_mem[6343];

	memory[1586][0] = temp_mem[6344];
	memory[1586][1] = temp_mem[6345];
	memory[1586][2] = temp_mem[6346];
	memory[1586][3] = temp_mem[6347];

	memory[1587][0] = temp_mem[6348];
	memory[1587][1] = temp_mem[6349];
	memory[1587][2] = temp_mem[6350];
	memory[1587][3] = temp_mem[6351];

	memory[1588][0] = temp_mem[6352];
	memory[1588][1] = temp_mem[6353];
	memory[1588][2] = temp_mem[6354];
	memory[1588][3] = temp_mem[6355];

	memory[1589][0] = temp_mem[6356];
	memory[1589][1] = temp_mem[6357];
	memory[1589][2] = temp_mem[6358];
	memory[1589][3] = temp_mem[6359];

	memory[1590][0] = temp_mem[6360];
	memory[1590][1] = temp_mem[6361];
	memory[1590][2] = temp_mem[6362];
	memory[1590][3] = temp_mem[6363];

	memory[1591][0] = temp_mem[6364];
	memory[1591][1] = temp_mem[6365];
	memory[1591][2] = temp_mem[6366];
	memory[1591][3] = temp_mem[6367];

	memory[1592][0] = temp_mem[6368];
	memory[1592][1] = temp_mem[6369];
	memory[1592][2] = temp_mem[6370];
	memory[1592][3] = temp_mem[6371];

	memory[1593][0] = temp_mem[6372];
	memory[1593][1] = temp_mem[6373];
	memory[1593][2] = temp_mem[6374];
	memory[1593][3] = temp_mem[6375];

	memory[1594][0] = temp_mem[6376];
	memory[1594][1] = temp_mem[6377];
	memory[1594][2] = temp_mem[6378];
	memory[1594][3] = temp_mem[6379];

	memory[1595][0] = temp_mem[6380];
	memory[1595][1] = temp_mem[6381];
	memory[1595][2] = temp_mem[6382];
	memory[1595][3] = temp_mem[6383];

	memory[1596][0] = temp_mem[6384];
	memory[1596][1] = temp_mem[6385];
	memory[1596][2] = temp_mem[6386];
	memory[1596][3] = temp_mem[6387];

	memory[1597][0] = temp_mem[6388];
	memory[1597][1] = temp_mem[6389];
	memory[1597][2] = temp_mem[6390];
	memory[1597][3] = temp_mem[6391];

	memory[1598][0] = temp_mem[6392];
	memory[1598][1] = temp_mem[6393];
	memory[1598][2] = temp_mem[6394];
	memory[1598][3] = temp_mem[6395];

	memory[1599][0] = temp_mem[6396];
	memory[1599][1] = temp_mem[6397];
	memory[1599][2] = temp_mem[6398];
	memory[1599][3] = temp_mem[6399];

	memory[1600][0] = temp_mem[6400];
	memory[1600][1] = temp_mem[6401];
	memory[1600][2] = temp_mem[6402];
	memory[1600][3] = temp_mem[6403];

	memory[1601][0] = temp_mem[6404];
	memory[1601][1] = temp_mem[6405];
	memory[1601][2] = temp_mem[6406];
	memory[1601][3] = temp_mem[6407];

	memory[1602][0] = temp_mem[6408];
	memory[1602][1] = temp_mem[6409];
	memory[1602][2] = temp_mem[6410];
	memory[1602][3] = temp_mem[6411];

	memory[1603][0] = temp_mem[6412];
	memory[1603][1] = temp_mem[6413];
	memory[1603][2] = temp_mem[6414];
	memory[1603][3] = temp_mem[6415];

	memory[1604][0] = temp_mem[6416];
	memory[1604][1] = temp_mem[6417];
	memory[1604][2] = temp_mem[6418];
	memory[1604][3] = temp_mem[6419];

	memory[1605][0] = temp_mem[6420];
	memory[1605][1] = temp_mem[6421];
	memory[1605][2] = temp_mem[6422];
	memory[1605][3] = temp_mem[6423];

	memory[1606][0] = temp_mem[6424];
	memory[1606][1] = temp_mem[6425];
	memory[1606][2] = temp_mem[6426];
	memory[1606][3] = temp_mem[6427];

	memory[1607][0] = temp_mem[6428];
	memory[1607][1] = temp_mem[6429];
	memory[1607][2] = temp_mem[6430];
	memory[1607][3] = temp_mem[6431];

	memory[1608][0] = temp_mem[6432];
	memory[1608][1] = temp_mem[6433];
	memory[1608][2] = temp_mem[6434];
	memory[1608][3] = temp_mem[6435];

	memory[1609][0] = temp_mem[6436];
	memory[1609][1] = temp_mem[6437];
	memory[1609][2] = temp_mem[6438];
	memory[1609][3] = temp_mem[6439];

	memory[1610][0] = temp_mem[6440];
	memory[1610][1] = temp_mem[6441];
	memory[1610][2] = temp_mem[6442];
	memory[1610][3] = temp_mem[6443];

	memory[1611][0] = temp_mem[6444];
	memory[1611][1] = temp_mem[6445];
	memory[1611][2] = temp_mem[6446];
	memory[1611][3] = temp_mem[6447];

	memory[1612][0] = temp_mem[6448];
	memory[1612][1] = temp_mem[6449];
	memory[1612][2] = temp_mem[6450];
	memory[1612][3] = temp_mem[6451];

	memory[1613][0] = temp_mem[6452];
	memory[1613][1] = temp_mem[6453];
	memory[1613][2] = temp_mem[6454];
	memory[1613][3] = temp_mem[6455];

	memory[1614][0] = temp_mem[6456];
	memory[1614][1] = temp_mem[6457];
	memory[1614][2] = temp_mem[6458];
	memory[1614][3] = temp_mem[6459];

	memory[1615][0] = temp_mem[6460];
	memory[1615][1] = temp_mem[6461];
	memory[1615][2] = temp_mem[6462];
	memory[1615][3] = temp_mem[6463];

	memory[1616][0] = temp_mem[6464];
	memory[1616][1] = temp_mem[6465];
	memory[1616][2] = temp_mem[6466];
	memory[1616][3] = temp_mem[6467];

	memory[1617][0] = temp_mem[6468];
	memory[1617][1] = temp_mem[6469];
	memory[1617][2] = temp_mem[6470];
	memory[1617][3] = temp_mem[6471];

	memory[1618][0] = temp_mem[6472];
	memory[1618][1] = temp_mem[6473];
	memory[1618][2] = temp_mem[6474];
	memory[1618][3] = temp_mem[6475];

	memory[1619][0] = temp_mem[6476];
	memory[1619][1] = temp_mem[6477];
	memory[1619][2] = temp_mem[6478];
	memory[1619][3] = temp_mem[6479];

	memory[1620][0] = temp_mem[6480];
	memory[1620][1] = temp_mem[6481];
	memory[1620][2] = temp_mem[6482];
	memory[1620][3] = temp_mem[6483];

	memory[1621][0] = temp_mem[6484];
	memory[1621][1] = temp_mem[6485];
	memory[1621][2] = temp_mem[6486];
	memory[1621][3] = temp_mem[6487];

	memory[1622][0] = temp_mem[6488];
	memory[1622][1] = temp_mem[6489];
	memory[1622][2] = temp_mem[6490];
	memory[1622][3] = temp_mem[6491];

	memory[1623][0] = temp_mem[6492];
	memory[1623][1] = temp_mem[6493];
	memory[1623][2] = temp_mem[6494];
	memory[1623][3] = temp_mem[6495];

	memory[1624][0] = temp_mem[6496];
	memory[1624][1] = temp_mem[6497];
	memory[1624][2] = temp_mem[6498];
	memory[1624][3] = temp_mem[6499];

	memory[1625][0] = temp_mem[6500];
	memory[1625][1] = temp_mem[6501];
	memory[1625][2] = temp_mem[6502];
	memory[1625][3] = temp_mem[6503];

	memory[1626][0] = temp_mem[6504];
	memory[1626][1] = temp_mem[6505];
	memory[1626][2] = temp_mem[6506];
	memory[1626][3] = temp_mem[6507];

	memory[1627][0] = temp_mem[6508];
	memory[1627][1] = temp_mem[6509];
	memory[1627][2] = temp_mem[6510];
	memory[1627][3] = temp_mem[6511];

	memory[1628][0] = temp_mem[6512];
	memory[1628][1] = temp_mem[6513];
	memory[1628][2] = temp_mem[6514];
	memory[1628][3] = temp_mem[6515];

	memory[1629][0] = temp_mem[6516];
	memory[1629][1] = temp_mem[6517];
	memory[1629][2] = temp_mem[6518];
	memory[1629][3] = temp_mem[6519];

	memory[1630][0] = temp_mem[6520];
	memory[1630][1] = temp_mem[6521];
	memory[1630][2] = temp_mem[6522];
	memory[1630][3] = temp_mem[6523];

	memory[1631][0] = temp_mem[6524];
	memory[1631][1] = temp_mem[6525];
	memory[1631][2] = temp_mem[6526];
	memory[1631][3] = temp_mem[6527];

	memory[1632][0] = temp_mem[6528];
	memory[1632][1] = temp_mem[6529];
	memory[1632][2] = temp_mem[6530];
	memory[1632][3] = temp_mem[6531];

	memory[1633][0] = temp_mem[6532];
	memory[1633][1] = temp_mem[6533];
	memory[1633][2] = temp_mem[6534];
	memory[1633][3] = temp_mem[6535];

	memory[1634][0] = temp_mem[6536];
	memory[1634][1] = temp_mem[6537];
	memory[1634][2] = temp_mem[6538];
	memory[1634][3] = temp_mem[6539];

	memory[1635][0] = temp_mem[6540];
	memory[1635][1] = temp_mem[6541];
	memory[1635][2] = temp_mem[6542];
	memory[1635][3] = temp_mem[6543];

	memory[1636][0] = temp_mem[6544];
	memory[1636][1] = temp_mem[6545];
	memory[1636][2] = temp_mem[6546];
	memory[1636][3] = temp_mem[6547];

	memory[1637][0] = temp_mem[6548];
	memory[1637][1] = temp_mem[6549];
	memory[1637][2] = temp_mem[6550];
	memory[1637][3] = temp_mem[6551];

	memory[1638][0] = temp_mem[6552];
	memory[1638][1] = temp_mem[6553];
	memory[1638][2] = temp_mem[6554];
	memory[1638][3] = temp_mem[6555];

	memory[1639][0] = temp_mem[6556];
	memory[1639][1] = temp_mem[6557];
	memory[1639][2] = temp_mem[6558];
	memory[1639][3] = temp_mem[6559];

	memory[1640][0] = temp_mem[6560];
	memory[1640][1] = temp_mem[6561];
	memory[1640][2] = temp_mem[6562];
	memory[1640][3] = temp_mem[6563];

	memory[1641][0] = temp_mem[6564];
	memory[1641][1] = temp_mem[6565];
	memory[1641][2] = temp_mem[6566];
	memory[1641][3] = temp_mem[6567];

	memory[1642][0] = temp_mem[6568];
	memory[1642][1] = temp_mem[6569];
	memory[1642][2] = temp_mem[6570];
	memory[1642][3] = temp_mem[6571];

	memory[1643][0] = temp_mem[6572];
	memory[1643][1] = temp_mem[6573];
	memory[1643][2] = temp_mem[6574];
	memory[1643][3] = temp_mem[6575];

	memory[1644][0] = temp_mem[6576];
	memory[1644][1] = temp_mem[6577];
	memory[1644][2] = temp_mem[6578];
	memory[1644][3] = temp_mem[6579];

	memory[1645][0] = temp_mem[6580];
	memory[1645][1] = temp_mem[6581];
	memory[1645][2] = temp_mem[6582];
	memory[1645][3] = temp_mem[6583];

	memory[1646][0] = temp_mem[6584];
	memory[1646][1] = temp_mem[6585];
	memory[1646][2] = temp_mem[6586];
	memory[1646][3] = temp_mem[6587];

	memory[1647][0] = temp_mem[6588];
	memory[1647][1] = temp_mem[6589];
	memory[1647][2] = temp_mem[6590];
	memory[1647][3] = temp_mem[6591];

	memory[1648][0] = temp_mem[6592];
	memory[1648][1] = temp_mem[6593];
	memory[1648][2] = temp_mem[6594];
	memory[1648][3] = temp_mem[6595];

	memory[1649][0] = temp_mem[6596];
	memory[1649][1] = temp_mem[6597];
	memory[1649][2] = temp_mem[6598];
	memory[1649][3] = temp_mem[6599];

	memory[1650][0] = temp_mem[6600];
	memory[1650][1] = temp_mem[6601];
	memory[1650][2] = temp_mem[6602];
	memory[1650][3] = temp_mem[6603];

	memory[1651][0] = temp_mem[6604];
	memory[1651][1] = temp_mem[6605];
	memory[1651][2] = temp_mem[6606];
	memory[1651][3] = temp_mem[6607];

	memory[1652][0] = temp_mem[6608];
	memory[1652][1] = temp_mem[6609];
	memory[1652][2] = temp_mem[6610];
	memory[1652][3] = temp_mem[6611];

	memory[1653][0] = temp_mem[6612];
	memory[1653][1] = temp_mem[6613];
	memory[1653][2] = temp_mem[6614];
	memory[1653][3] = temp_mem[6615];

	memory[1654][0] = temp_mem[6616];
	memory[1654][1] = temp_mem[6617];
	memory[1654][2] = temp_mem[6618];
	memory[1654][3] = temp_mem[6619];

	memory[1655][0] = temp_mem[6620];
	memory[1655][1] = temp_mem[6621];
	memory[1655][2] = temp_mem[6622];
	memory[1655][3] = temp_mem[6623];

	memory[1656][0] = temp_mem[6624];
	memory[1656][1] = temp_mem[6625];
	memory[1656][2] = temp_mem[6626];
	memory[1656][3] = temp_mem[6627];

	memory[1657][0] = temp_mem[6628];
	memory[1657][1] = temp_mem[6629];
	memory[1657][2] = temp_mem[6630];
	memory[1657][3] = temp_mem[6631];

	memory[1658][0] = temp_mem[6632];
	memory[1658][1] = temp_mem[6633];
	memory[1658][2] = temp_mem[6634];
	memory[1658][3] = temp_mem[6635];

	memory[1659][0] = temp_mem[6636];
	memory[1659][1] = temp_mem[6637];
	memory[1659][2] = temp_mem[6638];
	memory[1659][3] = temp_mem[6639];

	memory[1660][0] = temp_mem[6640];
	memory[1660][1] = temp_mem[6641];
	memory[1660][2] = temp_mem[6642];
	memory[1660][3] = temp_mem[6643];

	memory[1661][0] = temp_mem[6644];
	memory[1661][1] = temp_mem[6645];
	memory[1661][2] = temp_mem[6646];
	memory[1661][3] = temp_mem[6647];

	memory[1662][0] = temp_mem[6648];
	memory[1662][1] = temp_mem[6649];
	memory[1662][2] = temp_mem[6650];
	memory[1662][3] = temp_mem[6651];

	memory[1663][0] = temp_mem[6652];
	memory[1663][1] = temp_mem[6653];
	memory[1663][2] = temp_mem[6654];
	memory[1663][3] = temp_mem[6655];

	memory[1664][0] = temp_mem[6656];
	memory[1664][1] = temp_mem[6657];
	memory[1664][2] = temp_mem[6658];
	memory[1664][3] = temp_mem[6659];

	memory[1665][0] = temp_mem[6660];
	memory[1665][1] = temp_mem[6661];
	memory[1665][2] = temp_mem[6662];
	memory[1665][3] = temp_mem[6663];

	memory[1666][0] = temp_mem[6664];
	memory[1666][1] = temp_mem[6665];
	memory[1666][2] = temp_mem[6666];
	memory[1666][3] = temp_mem[6667];

	memory[1667][0] = temp_mem[6668];
	memory[1667][1] = temp_mem[6669];
	memory[1667][2] = temp_mem[6670];
	memory[1667][3] = temp_mem[6671];

	memory[1668][0] = temp_mem[6672];
	memory[1668][1] = temp_mem[6673];
	memory[1668][2] = temp_mem[6674];
	memory[1668][3] = temp_mem[6675];

	memory[1669][0] = temp_mem[6676];
	memory[1669][1] = temp_mem[6677];
	memory[1669][2] = temp_mem[6678];
	memory[1669][3] = temp_mem[6679];

	memory[1670][0] = temp_mem[6680];
	memory[1670][1] = temp_mem[6681];
	memory[1670][2] = temp_mem[6682];
	memory[1670][3] = temp_mem[6683];

	memory[1671][0] = temp_mem[6684];
	memory[1671][1] = temp_mem[6685];
	memory[1671][2] = temp_mem[6686];
	memory[1671][3] = temp_mem[6687];

	memory[1672][0] = temp_mem[6688];
	memory[1672][1] = temp_mem[6689];
	memory[1672][2] = temp_mem[6690];
	memory[1672][3] = temp_mem[6691];

	memory[1673][0] = temp_mem[6692];
	memory[1673][1] = temp_mem[6693];
	memory[1673][2] = temp_mem[6694];
	memory[1673][3] = temp_mem[6695];

	memory[1674][0] = temp_mem[6696];
	memory[1674][1] = temp_mem[6697];
	memory[1674][2] = temp_mem[6698];
	memory[1674][3] = temp_mem[6699];

	memory[1675][0] = temp_mem[6700];
	memory[1675][1] = temp_mem[6701];
	memory[1675][2] = temp_mem[6702];
	memory[1675][3] = temp_mem[6703];

	memory[1676][0] = temp_mem[6704];
	memory[1676][1] = temp_mem[6705];
	memory[1676][2] = temp_mem[6706];
	memory[1676][3] = temp_mem[6707];

	memory[1677][0] = temp_mem[6708];
	memory[1677][1] = temp_mem[6709];
	memory[1677][2] = temp_mem[6710];
	memory[1677][3] = temp_mem[6711];

	memory[1678][0] = temp_mem[6712];
	memory[1678][1] = temp_mem[6713];
	memory[1678][2] = temp_mem[6714];
	memory[1678][3] = temp_mem[6715];

	memory[1679][0] = temp_mem[6716];
	memory[1679][1] = temp_mem[6717];
	memory[1679][2] = temp_mem[6718];
	memory[1679][3] = temp_mem[6719];

	memory[1680][0] = temp_mem[6720];
	memory[1680][1] = temp_mem[6721];
	memory[1680][2] = temp_mem[6722];
	memory[1680][3] = temp_mem[6723];

	memory[1681][0] = temp_mem[6724];
	memory[1681][1] = temp_mem[6725];
	memory[1681][2] = temp_mem[6726];
	memory[1681][3] = temp_mem[6727];

	memory[1682][0] = temp_mem[6728];
	memory[1682][1] = temp_mem[6729];
	memory[1682][2] = temp_mem[6730];
	memory[1682][3] = temp_mem[6731];

	memory[1683][0] = temp_mem[6732];
	memory[1683][1] = temp_mem[6733];
	memory[1683][2] = temp_mem[6734];
	memory[1683][3] = temp_mem[6735];

	memory[1684][0] = temp_mem[6736];
	memory[1684][1] = temp_mem[6737];
	memory[1684][2] = temp_mem[6738];
	memory[1684][3] = temp_mem[6739];

	memory[1685][0] = temp_mem[6740];
	memory[1685][1] = temp_mem[6741];
	memory[1685][2] = temp_mem[6742];
	memory[1685][3] = temp_mem[6743];

	memory[1686][0] = temp_mem[6744];
	memory[1686][1] = temp_mem[6745];
	memory[1686][2] = temp_mem[6746];
	memory[1686][3] = temp_mem[6747];

	memory[1687][0] = temp_mem[6748];
	memory[1687][1] = temp_mem[6749];
	memory[1687][2] = temp_mem[6750];
	memory[1687][3] = temp_mem[6751];

	memory[1688][0] = temp_mem[6752];
	memory[1688][1] = temp_mem[6753];
	memory[1688][2] = temp_mem[6754];
	memory[1688][3] = temp_mem[6755];

	memory[1689][0] = temp_mem[6756];
	memory[1689][1] = temp_mem[6757];
	memory[1689][2] = temp_mem[6758];
	memory[1689][3] = temp_mem[6759];

	memory[1690][0] = temp_mem[6760];
	memory[1690][1] = temp_mem[6761];
	memory[1690][2] = temp_mem[6762];
	memory[1690][3] = temp_mem[6763];

	memory[1691][0] = temp_mem[6764];
	memory[1691][1] = temp_mem[6765];
	memory[1691][2] = temp_mem[6766];
	memory[1691][3] = temp_mem[6767];

	memory[1692][0] = temp_mem[6768];
	memory[1692][1] = temp_mem[6769];
	memory[1692][2] = temp_mem[6770];
	memory[1692][3] = temp_mem[6771];

	memory[1693][0] = temp_mem[6772];
	memory[1693][1] = temp_mem[6773];
	memory[1693][2] = temp_mem[6774];
	memory[1693][3] = temp_mem[6775];

	memory[1694][0] = temp_mem[6776];
	memory[1694][1] = temp_mem[6777];
	memory[1694][2] = temp_mem[6778];
	memory[1694][3] = temp_mem[6779];

	memory[1695][0] = temp_mem[6780];
	memory[1695][1] = temp_mem[6781];
	memory[1695][2] = temp_mem[6782];
	memory[1695][3] = temp_mem[6783];

	memory[1696][0] = temp_mem[6784];
	memory[1696][1] = temp_mem[6785];
	memory[1696][2] = temp_mem[6786];
	memory[1696][3] = temp_mem[6787];

	memory[1697][0] = temp_mem[6788];
	memory[1697][1] = temp_mem[6789];
	memory[1697][2] = temp_mem[6790];
	memory[1697][3] = temp_mem[6791];

	memory[1698][0] = temp_mem[6792];
	memory[1698][1] = temp_mem[6793];
	memory[1698][2] = temp_mem[6794];
	memory[1698][3] = temp_mem[6795];

	memory[1699][0] = temp_mem[6796];
	memory[1699][1] = temp_mem[6797];
	memory[1699][2] = temp_mem[6798];
	memory[1699][3] = temp_mem[6799];

	memory[1700][0] = temp_mem[6800];
	memory[1700][1] = temp_mem[6801];
	memory[1700][2] = temp_mem[6802];
	memory[1700][3] = temp_mem[6803];

	memory[1701][0] = temp_mem[6804];
	memory[1701][1] = temp_mem[6805];
	memory[1701][2] = temp_mem[6806];
	memory[1701][3] = temp_mem[6807];

	memory[1702][0] = temp_mem[6808];
	memory[1702][1] = temp_mem[6809];
	memory[1702][2] = temp_mem[6810];
	memory[1702][3] = temp_mem[6811];

	memory[1703][0] = temp_mem[6812];
	memory[1703][1] = temp_mem[6813];
	memory[1703][2] = temp_mem[6814];
	memory[1703][3] = temp_mem[6815];

	memory[1704][0] = temp_mem[6816];
	memory[1704][1] = temp_mem[6817];
	memory[1704][2] = temp_mem[6818];
	memory[1704][3] = temp_mem[6819];

	memory[1705][0] = temp_mem[6820];
	memory[1705][1] = temp_mem[6821];
	memory[1705][2] = temp_mem[6822];
	memory[1705][3] = temp_mem[6823];

	memory[1706][0] = temp_mem[6824];
	memory[1706][1] = temp_mem[6825];
	memory[1706][2] = temp_mem[6826];
	memory[1706][3] = temp_mem[6827];

	memory[1707][0] = temp_mem[6828];
	memory[1707][1] = temp_mem[6829];
	memory[1707][2] = temp_mem[6830];
	memory[1707][3] = temp_mem[6831];

	memory[1708][0] = temp_mem[6832];
	memory[1708][1] = temp_mem[6833];
	memory[1708][2] = temp_mem[6834];
	memory[1708][3] = temp_mem[6835];

	memory[1709][0] = temp_mem[6836];
	memory[1709][1] = temp_mem[6837];
	memory[1709][2] = temp_mem[6838];
	memory[1709][3] = temp_mem[6839];

	memory[1710][0] = temp_mem[6840];
	memory[1710][1] = temp_mem[6841];
	memory[1710][2] = temp_mem[6842];
	memory[1710][3] = temp_mem[6843];

	memory[1711][0] = temp_mem[6844];
	memory[1711][1] = temp_mem[6845];
	memory[1711][2] = temp_mem[6846];
	memory[1711][3] = temp_mem[6847];

	memory[1712][0] = temp_mem[6848];
	memory[1712][1] = temp_mem[6849];
	memory[1712][2] = temp_mem[6850];
	memory[1712][3] = temp_mem[6851];

	memory[1713][0] = temp_mem[6852];
	memory[1713][1] = temp_mem[6853];
	memory[1713][2] = temp_mem[6854];
	memory[1713][3] = temp_mem[6855];

	memory[1714][0] = temp_mem[6856];
	memory[1714][1] = temp_mem[6857];
	memory[1714][2] = temp_mem[6858];
	memory[1714][3] = temp_mem[6859];

	memory[1715][0] = temp_mem[6860];
	memory[1715][1] = temp_mem[6861];
	memory[1715][2] = temp_mem[6862];
	memory[1715][3] = temp_mem[6863];

	memory[1716][0] = temp_mem[6864];
	memory[1716][1] = temp_mem[6865];
	memory[1716][2] = temp_mem[6866];
	memory[1716][3] = temp_mem[6867];

	memory[1717][0] = temp_mem[6868];
	memory[1717][1] = temp_mem[6869];
	memory[1717][2] = temp_mem[6870];
	memory[1717][3] = temp_mem[6871];

	memory[1718][0] = temp_mem[6872];
	memory[1718][1] = temp_mem[6873];
	memory[1718][2] = temp_mem[6874];
	memory[1718][3] = temp_mem[6875];

	memory[1719][0] = temp_mem[6876];
	memory[1719][1] = temp_mem[6877];
	memory[1719][2] = temp_mem[6878];
	memory[1719][3] = temp_mem[6879];

	memory[1720][0] = temp_mem[6880];
	memory[1720][1] = temp_mem[6881];
	memory[1720][2] = temp_mem[6882];
	memory[1720][3] = temp_mem[6883];

	memory[1721][0] = temp_mem[6884];
	memory[1721][1] = temp_mem[6885];
	memory[1721][2] = temp_mem[6886];
	memory[1721][3] = temp_mem[6887];

	memory[1722][0] = temp_mem[6888];
	memory[1722][1] = temp_mem[6889];
	memory[1722][2] = temp_mem[6890];
	memory[1722][3] = temp_mem[6891];

	memory[1723][0] = temp_mem[6892];
	memory[1723][1] = temp_mem[6893];
	memory[1723][2] = temp_mem[6894];
	memory[1723][3] = temp_mem[6895];

	memory[1724][0] = temp_mem[6896];
	memory[1724][1] = temp_mem[6897];
	memory[1724][2] = temp_mem[6898];
	memory[1724][3] = temp_mem[6899];

	memory[1725][0] = temp_mem[6900];
	memory[1725][1] = temp_mem[6901];
	memory[1725][2] = temp_mem[6902];
	memory[1725][3] = temp_mem[6903];

	memory[1726][0] = temp_mem[6904];
	memory[1726][1] = temp_mem[6905];
	memory[1726][2] = temp_mem[6906];
	memory[1726][3] = temp_mem[6907];

	memory[1727][0] = temp_mem[6908];
	memory[1727][1] = temp_mem[6909];
	memory[1727][2] = temp_mem[6910];
	memory[1727][3] = temp_mem[6911];

	memory[1728][0] = temp_mem[6912];
	memory[1728][1] = temp_mem[6913];
	memory[1728][2] = temp_mem[6914];
	memory[1728][3] = temp_mem[6915];

	memory[1729][0] = temp_mem[6916];
	memory[1729][1] = temp_mem[6917];
	memory[1729][2] = temp_mem[6918];
	memory[1729][3] = temp_mem[6919];

	memory[1730][0] = temp_mem[6920];
	memory[1730][1] = temp_mem[6921];
	memory[1730][2] = temp_mem[6922];
	memory[1730][3] = temp_mem[6923];

	memory[1731][0] = temp_mem[6924];
	memory[1731][1] = temp_mem[6925];
	memory[1731][2] = temp_mem[6926];
	memory[1731][3] = temp_mem[6927];

	memory[1732][0] = temp_mem[6928];
	memory[1732][1] = temp_mem[6929];
	memory[1732][2] = temp_mem[6930];
	memory[1732][3] = temp_mem[6931];

	memory[1733][0] = temp_mem[6932];
	memory[1733][1] = temp_mem[6933];
	memory[1733][2] = temp_mem[6934];
	memory[1733][3] = temp_mem[6935];

	memory[1734][0] = temp_mem[6936];
	memory[1734][1] = temp_mem[6937];
	memory[1734][2] = temp_mem[6938];
	memory[1734][3] = temp_mem[6939];

	memory[1735][0] = temp_mem[6940];
	memory[1735][1] = temp_mem[6941];
	memory[1735][2] = temp_mem[6942];
	memory[1735][3] = temp_mem[6943];

	memory[1736][0] = temp_mem[6944];
	memory[1736][1] = temp_mem[6945];
	memory[1736][2] = temp_mem[6946];
	memory[1736][3] = temp_mem[6947];

	memory[1737][0] = temp_mem[6948];
	memory[1737][1] = temp_mem[6949];
	memory[1737][2] = temp_mem[6950];
	memory[1737][3] = temp_mem[6951];

	memory[1738][0] = temp_mem[6952];
	memory[1738][1] = temp_mem[6953];
	memory[1738][2] = temp_mem[6954];
	memory[1738][3] = temp_mem[6955];

	memory[1739][0] = temp_mem[6956];
	memory[1739][1] = temp_mem[6957];
	memory[1739][2] = temp_mem[6958];
	memory[1739][3] = temp_mem[6959];

	memory[1740][0] = temp_mem[6960];
	memory[1740][1] = temp_mem[6961];
	memory[1740][2] = temp_mem[6962];
	memory[1740][3] = temp_mem[6963];

	memory[1741][0] = temp_mem[6964];
	memory[1741][1] = temp_mem[6965];
	memory[1741][2] = temp_mem[6966];
	memory[1741][3] = temp_mem[6967];

	memory[1742][0] = temp_mem[6968];
	memory[1742][1] = temp_mem[6969];
	memory[1742][2] = temp_mem[6970];
	memory[1742][3] = temp_mem[6971];

	memory[1743][0] = temp_mem[6972];
	memory[1743][1] = temp_mem[6973];
	memory[1743][2] = temp_mem[6974];
	memory[1743][3] = temp_mem[6975];

	memory[1744][0] = temp_mem[6976];
	memory[1744][1] = temp_mem[6977];
	memory[1744][2] = temp_mem[6978];
	memory[1744][3] = temp_mem[6979];

	memory[1745][0] = temp_mem[6980];
	memory[1745][1] = temp_mem[6981];
	memory[1745][2] = temp_mem[6982];
	memory[1745][3] = temp_mem[6983];

	memory[1746][0] = temp_mem[6984];
	memory[1746][1] = temp_mem[6985];
	memory[1746][2] = temp_mem[6986];
	memory[1746][3] = temp_mem[6987];

	memory[1747][0] = temp_mem[6988];
	memory[1747][1] = temp_mem[6989];
	memory[1747][2] = temp_mem[6990];
	memory[1747][3] = temp_mem[6991];

	memory[1748][0] = temp_mem[6992];
	memory[1748][1] = temp_mem[6993];
	memory[1748][2] = temp_mem[6994];
	memory[1748][3] = temp_mem[6995];

	memory[1749][0] = temp_mem[6996];
	memory[1749][1] = temp_mem[6997];
	memory[1749][2] = temp_mem[6998];
	memory[1749][3] = temp_mem[6999];

	memory[1750][0] = temp_mem[7000];
	memory[1750][1] = temp_mem[7001];
	memory[1750][2] = temp_mem[7002];
	memory[1750][3] = temp_mem[7003];

	memory[1751][0] = temp_mem[7004];
	memory[1751][1] = temp_mem[7005];
	memory[1751][2] = temp_mem[7006];
	memory[1751][3] = temp_mem[7007];

	memory[1752][0] = temp_mem[7008];
	memory[1752][1] = temp_mem[7009];
	memory[1752][2] = temp_mem[7010];
	memory[1752][3] = temp_mem[7011];

	memory[1753][0] = temp_mem[7012];
	memory[1753][1] = temp_mem[7013];
	memory[1753][2] = temp_mem[7014];
	memory[1753][3] = temp_mem[7015];

	memory[1754][0] = temp_mem[7016];
	memory[1754][1] = temp_mem[7017];
	memory[1754][2] = temp_mem[7018];
	memory[1754][3] = temp_mem[7019];

	memory[1755][0] = temp_mem[7020];
	memory[1755][1] = temp_mem[7021];
	memory[1755][2] = temp_mem[7022];
	memory[1755][3] = temp_mem[7023];

	memory[1756][0] = temp_mem[7024];
	memory[1756][1] = temp_mem[7025];
	memory[1756][2] = temp_mem[7026];
	memory[1756][3] = temp_mem[7027];

	memory[1757][0] = temp_mem[7028];
	memory[1757][1] = temp_mem[7029];
	memory[1757][2] = temp_mem[7030];
	memory[1757][3] = temp_mem[7031];

	memory[1758][0] = temp_mem[7032];
	memory[1758][1] = temp_mem[7033];
	memory[1758][2] = temp_mem[7034];
	memory[1758][3] = temp_mem[7035];

	memory[1759][0] = temp_mem[7036];
	memory[1759][1] = temp_mem[7037];
	memory[1759][2] = temp_mem[7038];
	memory[1759][3] = temp_mem[7039];

	memory[1760][0] = temp_mem[7040];
	memory[1760][1] = temp_mem[7041];
	memory[1760][2] = temp_mem[7042];
	memory[1760][3] = temp_mem[7043];

	memory[1761][0] = temp_mem[7044];
	memory[1761][1] = temp_mem[7045];
	memory[1761][2] = temp_mem[7046];
	memory[1761][3] = temp_mem[7047];

	memory[1762][0] = temp_mem[7048];
	memory[1762][1] = temp_mem[7049];
	memory[1762][2] = temp_mem[7050];
	memory[1762][3] = temp_mem[7051];

	memory[1763][0] = temp_mem[7052];
	memory[1763][1] = temp_mem[7053];
	memory[1763][2] = temp_mem[7054];
	memory[1763][3] = temp_mem[7055];

	memory[1764][0] = temp_mem[7056];
	memory[1764][1] = temp_mem[7057];
	memory[1764][2] = temp_mem[7058];
	memory[1764][3] = temp_mem[7059];

	memory[1765][0] = temp_mem[7060];
	memory[1765][1] = temp_mem[7061];
	memory[1765][2] = temp_mem[7062];
	memory[1765][3] = temp_mem[7063];

	memory[1766][0] = temp_mem[7064];
	memory[1766][1] = temp_mem[7065];
	memory[1766][2] = temp_mem[7066];
	memory[1766][3] = temp_mem[7067];

	memory[1767][0] = temp_mem[7068];
	memory[1767][1] = temp_mem[7069];
	memory[1767][2] = temp_mem[7070];
	memory[1767][3] = temp_mem[7071];

	memory[1768][0] = temp_mem[7072];
	memory[1768][1] = temp_mem[7073];
	memory[1768][2] = temp_mem[7074];
	memory[1768][3] = temp_mem[7075];

	memory[1769][0] = temp_mem[7076];
	memory[1769][1] = temp_mem[7077];
	memory[1769][2] = temp_mem[7078];
	memory[1769][3] = temp_mem[7079];

	memory[1770][0] = temp_mem[7080];
	memory[1770][1] = temp_mem[7081];
	memory[1770][2] = temp_mem[7082];
	memory[1770][3] = temp_mem[7083];

	memory[1771][0] = temp_mem[7084];
	memory[1771][1] = temp_mem[7085];
	memory[1771][2] = temp_mem[7086];
	memory[1771][3] = temp_mem[7087];

	memory[1772][0] = temp_mem[7088];
	memory[1772][1] = temp_mem[7089];
	memory[1772][2] = temp_mem[7090];
	memory[1772][3] = temp_mem[7091];

	memory[1773][0] = temp_mem[7092];
	memory[1773][1] = temp_mem[7093];
	memory[1773][2] = temp_mem[7094];
	memory[1773][3] = temp_mem[7095];

	memory[1774][0] = temp_mem[7096];
	memory[1774][1] = temp_mem[7097];
	memory[1774][2] = temp_mem[7098];
	memory[1774][3] = temp_mem[7099];

	memory[1775][0] = temp_mem[7100];
	memory[1775][1] = temp_mem[7101];
	memory[1775][2] = temp_mem[7102];
	memory[1775][3] = temp_mem[7103];

	memory[1776][0] = temp_mem[7104];
	memory[1776][1] = temp_mem[7105];
	memory[1776][2] = temp_mem[7106];
	memory[1776][3] = temp_mem[7107];

	memory[1777][0] = temp_mem[7108];
	memory[1777][1] = temp_mem[7109];
	memory[1777][2] = temp_mem[7110];
	memory[1777][3] = temp_mem[7111];

	memory[1778][0] = temp_mem[7112];
	memory[1778][1] = temp_mem[7113];
	memory[1778][2] = temp_mem[7114];
	memory[1778][3] = temp_mem[7115];

	memory[1779][0] = temp_mem[7116];
	memory[1779][1] = temp_mem[7117];
	memory[1779][2] = temp_mem[7118];
	memory[1779][3] = temp_mem[7119];

	memory[1780][0] = temp_mem[7120];
	memory[1780][1] = temp_mem[7121];
	memory[1780][2] = temp_mem[7122];
	memory[1780][3] = temp_mem[7123];

	memory[1781][0] = temp_mem[7124];
	memory[1781][1] = temp_mem[7125];
	memory[1781][2] = temp_mem[7126];
	memory[1781][3] = temp_mem[7127];

	memory[1782][0] = temp_mem[7128];
	memory[1782][1] = temp_mem[7129];
	memory[1782][2] = temp_mem[7130];
	memory[1782][3] = temp_mem[7131];

	memory[1783][0] = temp_mem[7132];
	memory[1783][1] = temp_mem[7133];
	memory[1783][2] = temp_mem[7134];
	memory[1783][3] = temp_mem[7135];

	memory[1784][0] = temp_mem[7136];
	memory[1784][1] = temp_mem[7137];
	memory[1784][2] = temp_mem[7138];
	memory[1784][3] = temp_mem[7139];

	memory[1785][0] = temp_mem[7140];
	memory[1785][1] = temp_mem[7141];
	memory[1785][2] = temp_mem[7142];
	memory[1785][3] = temp_mem[7143];

	memory[1786][0] = temp_mem[7144];
	memory[1786][1] = temp_mem[7145];
	memory[1786][2] = temp_mem[7146];
	memory[1786][3] = temp_mem[7147];

	memory[1787][0] = temp_mem[7148];
	memory[1787][1] = temp_mem[7149];
	memory[1787][2] = temp_mem[7150];
	memory[1787][3] = temp_mem[7151];

	memory[1788][0] = temp_mem[7152];
	memory[1788][1] = temp_mem[7153];
	memory[1788][2] = temp_mem[7154];
	memory[1788][3] = temp_mem[7155];

	memory[1789][0] = temp_mem[7156];
	memory[1789][1] = temp_mem[7157];
	memory[1789][2] = temp_mem[7158];
	memory[1789][3] = temp_mem[7159];

	memory[1790][0] = temp_mem[7160];
	memory[1790][1] = temp_mem[7161];
	memory[1790][2] = temp_mem[7162];
	memory[1790][3] = temp_mem[7163];

	memory[1791][0] = temp_mem[7164];
	memory[1791][1] = temp_mem[7165];
	memory[1791][2] = temp_mem[7166];
	memory[1791][3] = temp_mem[7167];

	memory[1792][0] = temp_mem[7168];
	memory[1792][1] = temp_mem[7169];
	memory[1792][2] = temp_mem[7170];
	memory[1792][3] = temp_mem[7171];

	memory[1793][0] = temp_mem[7172];
	memory[1793][1] = temp_mem[7173];
	memory[1793][2] = temp_mem[7174];
	memory[1793][3] = temp_mem[7175];

	memory[1794][0] = temp_mem[7176];
	memory[1794][1] = temp_mem[7177];
	memory[1794][2] = temp_mem[7178];
	memory[1794][3] = temp_mem[7179];

	memory[1795][0] = temp_mem[7180];
	memory[1795][1] = temp_mem[7181];
	memory[1795][2] = temp_mem[7182];
	memory[1795][3] = temp_mem[7183];

	memory[1796][0] = temp_mem[7184];
	memory[1796][1] = temp_mem[7185];
	memory[1796][2] = temp_mem[7186];
	memory[1796][3] = temp_mem[7187];

	memory[1797][0] = temp_mem[7188];
	memory[1797][1] = temp_mem[7189];
	memory[1797][2] = temp_mem[7190];
	memory[1797][3] = temp_mem[7191];

	memory[1798][0] = temp_mem[7192];
	memory[1798][1] = temp_mem[7193];
	memory[1798][2] = temp_mem[7194];
	memory[1798][3] = temp_mem[7195];

	memory[1799][0] = temp_mem[7196];
	memory[1799][1] = temp_mem[7197];
	memory[1799][2] = temp_mem[7198];
	memory[1799][3] = temp_mem[7199];

	memory[1800][0] = temp_mem[7200];
	memory[1800][1] = temp_mem[7201];
	memory[1800][2] = temp_mem[7202];
	memory[1800][3] = temp_mem[7203];

	memory[1801][0] = temp_mem[7204];
	memory[1801][1] = temp_mem[7205];
	memory[1801][2] = temp_mem[7206];
	memory[1801][3] = temp_mem[7207];

	memory[1802][0] = temp_mem[7208];
	memory[1802][1] = temp_mem[7209];
	memory[1802][2] = temp_mem[7210];
	memory[1802][3] = temp_mem[7211];

	memory[1803][0] = temp_mem[7212];
	memory[1803][1] = temp_mem[7213];
	memory[1803][2] = temp_mem[7214];
	memory[1803][3] = temp_mem[7215];

	memory[1804][0] = temp_mem[7216];
	memory[1804][1] = temp_mem[7217];
	memory[1804][2] = temp_mem[7218];
	memory[1804][3] = temp_mem[7219];

	memory[1805][0] = temp_mem[7220];
	memory[1805][1] = temp_mem[7221];
	memory[1805][2] = temp_mem[7222];
	memory[1805][3] = temp_mem[7223];

	memory[1806][0] = temp_mem[7224];
	memory[1806][1] = temp_mem[7225];
	memory[1806][2] = temp_mem[7226];
	memory[1806][3] = temp_mem[7227];

	memory[1807][0] = temp_mem[7228];
	memory[1807][1] = temp_mem[7229];
	memory[1807][2] = temp_mem[7230];
	memory[1807][3] = temp_mem[7231];

	memory[1808][0] = temp_mem[7232];
	memory[1808][1] = temp_mem[7233];
	memory[1808][2] = temp_mem[7234];
	memory[1808][3] = temp_mem[7235];

	memory[1809][0] = temp_mem[7236];
	memory[1809][1] = temp_mem[7237];
	memory[1809][2] = temp_mem[7238];
	memory[1809][3] = temp_mem[7239];

	memory[1810][0] = temp_mem[7240];
	memory[1810][1] = temp_mem[7241];
	memory[1810][2] = temp_mem[7242];
	memory[1810][3] = temp_mem[7243];

	memory[1811][0] = temp_mem[7244];
	memory[1811][1] = temp_mem[7245];
	memory[1811][2] = temp_mem[7246];
	memory[1811][3] = temp_mem[7247];

	memory[1812][0] = temp_mem[7248];
	memory[1812][1] = temp_mem[7249];
	memory[1812][2] = temp_mem[7250];
	memory[1812][3] = temp_mem[7251];

	memory[1813][0] = temp_mem[7252];
	memory[1813][1] = temp_mem[7253];
	memory[1813][2] = temp_mem[7254];
	memory[1813][3] = temp_mem[7255];

	memory[1814][0] = temp_mem[7256];
	memory[1814][1] = temp_mem[7257];
	memory[1814][2] = temp_mem[7258];
	memory[1814][3] = temp_mem[7259];

	memory[1815][0] = temp_mem[7260];
	memory[1815][1] = temp_mem[7261];
	memory[1815][2] = temp_mem[7262];
	memory[1815][3] = temp_mem[7263];

	memory[1816][0] = temp_mem[7264];
	memory[1816][1] = temp_mem[7265];
	memory[1816][2] = temp_mem[7266];
	memory[1816][3] = temp_mem[7267];

	memory[1817][0] = temp_mem[7268];
	memory[1817][1] = temp_mem[7269];
	memory[1817][2] = temp_mem[7270];
	memory[1817][3] = temp_mem[7271];

	memory[1818][0] = temp_mem[7272];
	memory[1818][1] = temp_mem[7273];
	memory[1818][2] = temp_mem[7274];
	memory[1818][3] = temp_mem[7275];

	memory[1819][0] = temp_mem[7276];
	memory[1819][1] = temp_mem[7277];
	memory[1819][2] = temp_mem[7278];
	memory[1819][3] = temp_mem[7279];

	memory[1820][0] = temp_mem[7280];
	memory[1820][1] = temp_mem[7281];
	memory[1820][2] = temp_mem[7282];
	memory[1820][3] = temp_mem[7283];

	memory[1821][0] = temp_mem[7284];
	memory[1821][1] = temp_mem[7285];
	memory[1821][2] = temp_mem[7286];
	memory[1821][3] = temp_mem[7287];

	memory[1822][0] = temp_mem[7288];
	memory[1822][1] = temp_mem[7289];
	memory[1822][2] = temp_mem[7290];
	memory[1822][3] = temp_mem[7291];

	memory[1823][0] = temp_mem[7292];
	memory[1823][1] = temp_mem[7293];
	memory[1823][2] = temp_mem[7294];
	memory[1823][3] = temp_mem[7295];

	memory[1824][0] = temp_mem[7296];
	memory[1824][1] = temp_mem[7297];
	memory[1824][2] = temp_mem[7298];
	memory[1824][3] = temp_mem[7299];

	memory[1825][0] = temp_mem[7300];
	memory[1825][1] = temp_mem[7301];
	memory[1825][2] = temp_mem[7302];
	memory[1825][3] = temp_mem[7303];

	memory[1826][0] = temp_mem[7304];
	memory[1826][1] = temp_mem[7305];
	memory[1826][2] = temp_mem[7306];
	memory[1826][3] = temp_mem[7307];

	memory[1827][0] = temp_mem[7308];
	memory[1827][1] = temp_mem[7309];
	memory[1827][2] = temp_mem[7310];
	memory[1827][3] = temp_mem[7311];

	memory[1828][0] = temp_mem[7312];
	memory[1828][1] = temp_mem[7313];
	memory[1828][2] = temp_mem[7314];
	memory[1828][3] = temp_mem[7315];

	memory[1829][0] = temp_mem[7316];
	memory[1829][1] = temp_mem[7317];
	memory[1829][2] = temp_mem[7318];
	memory[1829][3] = temp_mem[7319];

	memory[1830][0] = temp_mem[7320];
	memory[1830][1] = temp_mem[7321];
	memory[1830][2] = temp_mem[7322];
	memory[1830][3] = temp_mem[7323];

	memory[1831][0] = temp_mem[7324];
	memory[1831][1] = temp_mem[7325];
	memory[1831][2] = temp_mem[7326];
	memory[1831][3] = temp_mem[7327];

	memory[1832][0] = temp_mem[7328];
	memory[1832][1] = temp_mem[7329];
	memory[1832][2] = temp_mem[7330];
	memory[1832][3] = temp_mem[7331];

	memory[1833][0] = temp_mem[7332];
	memory[1833][1] = temp_mem[7333];
	memory[1833][2] = temp_mem[7334];
	memory[1833][3] = temp_mem[7335];

	memory[1834][0] = temp_mem[7336];
	memory[1834][1] = temp_mem[7337];
	memory[1834][2] = temp_mem[7338];
	memory[1834][3] = temp_mem[7339];

	memory[1835][0] = temp_mem[7340];
	memory[1835][1] = temp_mem[7341];
	memory[1835][2] = temp_mem[7342];
	memory[1835][3] = temp_mem[7343];

	memory[1836][0] = temp_mem[7344];
	memory[1836][1] = temp_mem[7345];
	memory[1836][2] = temp_mem[7346];
	memory[1836][3] = temp_mem[7347];

	memory[1837][0] = temp_mem[7348];
	memory[1837][1] = temp_mem[7349];
	memory[1837][2] = temp_mem[7350];
	memory[1837][3] = temp_mem[7351];

	memory[1838][0] = temp_mem[7352];
	memory[1838][1] = temp_mem[7353];
	memory[1838][2] = temp_mem[7354];
	memory[1838][3] = temp_mem[7355];

	memory[1839][0] = temp_mem[7356];
	memory[1839][1] = temp_mem[7357];
	memory[1839][2] = temp_mem[7358];
	memory[1839][3] = temp_mem[7359];

	memory[1840][0] = temp_mem[7360];
	memory[1840][1] = temp_mem[7361];
	memory[1840][2] = temp_mem[7362];
	memory[1840][3] = temp_mem[7363];

	memory[1841][0] = temp_mem[7364];
	memory[1841][1] = temp_mem[7365];
	memory[1841][2] = temp_mem[7366];
	memory[1841][3] = temp_mem[7367];

	memory[1842][0] = temp_mem[7368];
	memory[1842][1] = temp_mem[7369];
	memory[1842][2] = temp_mem[7370];
	memory[1842][3] = temp_mem[7371];

	memory[1843][0] = temp_mem[7372];
	memory[1843][1] = temp_mem[7373];
	memory[1843][2] = temp_mem[7374];
	memory[1843][3] = temp_mem[7375];

	memory[1844][0] = temp_mem[7376];
	memory[1844][1] = temp_mem[7377];
	memory[1844][2] = temp_mem[7378];
	memory[1844][3] = temp_mem[7379];

	memory[1845][0] = temp_mem[7380];
	memory[1845][1] = temp_mem[7381];
	memory[1845][2] = temp_mem[7382];
	memory[1845][3] = temp_mem[7383];

	memory[1846][0] = temp_mem[7384];
	memory[1846][1] = temp_mem[7385];
	memory[1846][2] = temp_mem[7386];
	memory[1846][3] = temp_mem[7387];

	memory[1847][0] = temp_mem[7388];
	memory[1847][1] = temp_mem[7389];
	memory[1847][2] = temp_mem[7390];
	memory[1847][3] = temp_mem[7391];

	memory[1848][0] = temp_mem[7392];
	memory[1848][1] = temp_mem[7393];
	memory[1848][2] = temp_mem[7394];
	memory[1848][3] = temp_mem[7395];

	memory[1849][0] = temp_mem[7396];
	memory[1849][1] = temp_mem[7397];
	memory[1849][2] = temp_mem[7398];
	memory[1849][3] = temp_mem[7399];

	memory[1850][0] = temp_mem[7400];
	memory[1850][1] = temp_mem[7401];
	memory[1850][2] = temp_mem[7402];
	memory[1850][3] = temp_mem[7403];

	memory[1851][0] = temp_mem[7404];
	memory[1851][1] = temp_mem[7405];
	memory[1851][2] = temp_mem[7406];
	memory[1851][3] = temp_mem[7407];

	memory[1852][0] = temp_mem[7408];
	memory[1852][1] = temp_mem[7409];
	memory[1852][2] = temp_mem[7410];
	memory[1852][3] = temp_mem[7411];

	memory[1853][0] = temp_mem[7412];
	memory[1853][1] = temp_mem[7413];
	memory[1853][2] = temp_mem[7414];
	memory[1853][3] = temp_mem[7415];

	memory[1854][0] = temp_mem[7416];
	memory[1854][1] = temp_mem[7417];
	memory[1854][2] = temp_mem[7418];
	memory[1854][3] = temp_mem[7419];

	memory[1855][0] = temp_mem[7420];
	memory[1855][1] = temp_mem[7421];
	memory[1855][2] = temp_mem[7422];
	memory[1855][3] = temp_mem[7423];

	memory[1856][0] = temp_mem[7424];
	memory[1856][1] = temp_mem[7425];
	memory[1856][2] = temp_mem[7426];
	memory[1856][3] = temp_mem[7427];

	memory[1857][0] = temp_mem[7428];
	memory[1857][1] = temp_mem[7429];
	memory[1857][2] = temp_mem[7430];
	memory[1857][3] = temp_mem[7431];

	memory[1858][0] = temp_mem[7432];
	memory[1858][1] = temp_mem[7433];
	memory[1858][2] = temp_mem[7434];
	memory[1858][3] = temp_mem[7435];

	memory[1859][0] = temp_mem[7436];
	memory[1859][1] = temp_mem[7437];
	memory[1859][2] = temp_mem[7438];
	memory[1859][3] = temp_mem[7439];

	memory[1860][0] = temp_mem[7440];
	memory[1860][1] = temp_mem[7441];
	memory[1860][2] = temp_mem[7442];
	memory[1860][3] = temp_mem[7443];

	memory[1861][0] = temp_mem[7444];
	memory[1861][1] = temp_mem[7445];
	memory[1861][2] = temp_mem[7446];
	memory[1861][3] = temp_mem[7447];

	memory[1862][0] = temp_mem[7448];
	memory[1862][1] = temp_mem[7449];
	memory[1862][2] = temp_mem[7450];
	memory[1862][3] = temp_mem[7451];

	memory[1863][0] = temp_mem[7452];
	memory[1863][1] = temp_mem[7453];
	memory[1863][2] = temp_mem[7454];
	memory[1863][3] = temp_mem[7455];

	memory[1864][0] = temp_mem[7456];
	memory[1864][1] = temp_mem[7457];
	memory[1864][2] = temp_mem[7458];
	memory[1864][3] = temp_mem[7459];

	memory[1865][0] = temp_mem[7460];
	memory[1865][1] = temp_mem[7461];
	memory[1865][2] = temp_mem[7462];
	memory[1865][3] = temp_mem[7463];

	memory[1866][0] = temp_mem[7464];
	memory[1866][1] = temp_mem[7465];
	memory[1866][2] = temp_mem[7466];
	memory[1866][3] = temp_mem[7467];

	memory[1867][0] = temp_mem[7468];
	memory[1867][1] = temp_mem[7469];
	memory[1867][2] = temp_mem[7470];
	memory[1867][3] = temp_mem[7471];

	memory[1868][0] = temp_mem[7472];
	memory[1868][1] = temp_mem[7473];
	memory[1868][2] = temp_mem[7474];
	memory[1868][3] = temp_mem[7475];

	memory[1869][0] = temp_mem[7476];
	memory[1869][1] = temp_mem[7477];
	memory[1869][2] = temp_mem[7478];
	memory[1869][3] = temp_mem[7479];

	memory[1870][0] = temp_mem[7480];
	memory[1870][1] = temp_mem[7481];
	memory[1870][2] = temp_mem[7482];
	memory[1870][3] = temp_mem[7483];

	memory[1871][0] = temp_mem[7484];
	memory[1871][1] = temp_mem[7485];
	memory[1871][2] = temp_mem[7486];
	memory[1871][3] = temp_mem[7487];

	memory[1872][0] = temp_mem[7488];
	memory[1872][1] = temp_mem[7489];
	memory[1872][2] = temp_mem[7490];
	memory[1872][3] = temp_mem[7491];

	memory[1873][0] = temp_mem[7492];
	memory[1873][1] = temp_mem[7493];
	memory[1873][2] = temp_mem[7494];
	memory[1873][3] = temp_mem[7495];

	memory[1874][0] = temp_mem[7496];
	memory[1874][1] = temp_mem[7497];
	memory[1874][2] = temp_mem[7498];
	memory[1874][3] = temp_mem[7499];

	memory[1875][0] = temp_mem[7500];
	memory[1875][1] = temp_mem[7501];
	memory[1875][2] = temp_mem[7502];
	memory[1875][3] = temp_mem[7503];

	memory[1876][0] = temp_mem[7504];
	memory[1876][1] = temp_mem[7505];
	memory[1876][2] = temp_mem[7506];
	memory[1876][3] = temp_mem[7507];

	memory[1877][0] = temp_mem[7508];
	memory[1877][1] = temp_mem[7509];
	memory[1877][2] = temp_mem[7510];
	memory[1877][3] = temp_mem[7511];

	memory[1878][0] = temp_mem[7512];
	memory[1878][1] = temp_mem[7513];
	memory[1878][2] = temp_mem[7514];
	memory[1878][3] = temp_mem[7515];

	memory[1879][0] = temp_mem[7516];
	memory[1879][1] = temp_mem[7517];
	memory[1879][2] = temp_mem[7518];
	memory[1879][3] = temp_mem[7519];

	memory[1880][0] = temp_mem[7520];
	memory[1880][1] = temp_mem[7521];
	memory[1880][2] = temp_mem[7522];
	memory[1880][3] = temp_mem[7523];

	memory[1881][0] = temp_mem[7524];
	memory[1881][1] = temp_mem[7525];
	memory[1881][2] = temp_mem[7526];
	memory[1881][3] = temp_mem[7527];

	memory[1882][0] = temp_mem[7528];
	memory[1882][1] = temp_mem[7529];
	memory[1882][2] = temp_mem[7530];
	memory[1882][3] = temp_mem[7531];

	memory[1883][0] = temp_mem[7532];
	memory[1883][1] = temp_mem[7533];
	memory[1883][2] = temp_mem[7534];
	memory[1883][3] = temp_mem[7535];

	memory[1884][0] = temp_mem[7536];
	memory[1884][1] = temp_mem[7537];
	memory[1884][2] = temp_mem[7538];
	memory[1884][3] = temp_mem[7539];

	memory[1885][0] = temp_mem[7540];
	memory[1885][1] = temp_mem[7541];
	memory[1885][2] = temp_mem[7542];
	memory[1885][3] = temp_mem[7543];

	memory[1886][0] = temp_mem[7544];
	memory[1886][1] = temp_mem[7545];
	memory[1886][2] = temp_mem[7546];
	memory[1886][3] = temp_mem[7547];

	memory[1887][0] = temp_mem[7548];
	memory[1887][1] = temp_mem[7549];
	memory[1887][2] = temp_mem[7550];
	memory[1887][3] = temp_mem[7551];

	memory[1888][0] = temp_mem[7552];
	memory[1888][1] = temp_mem[7553];
	memory[1888][2] = temp_mem[7554];
	memory[1888][3] = temp_mem[7555];

	memory[1889][0] = temp_mem[7556];
	memory[1889][1] = temp_mem[7557];
	memory[1889][2] = temp_mem[7558];
	memory[1889][3] = temp_mem[7559];

	memory[1890][0] = temp_mem[7560];
	memory[1890][1] = temp_mem[7561];
	memory[1890][2] = temp_mem[7562];
	memory[1890][3] = temp_mem[7563];

	memory[1891][0] = temp_mem[7564];
	memory[1891][1] = temp_mem[7565];
	memory[1891][2] = temp_mem[7566];
	memory[1891][3] = temp_mem[7567];

	memory[1892][0] = temp_mem[7568];
	memory[1892][1] = temp_mem[7569];
	memory[1892][2] = temp_mem[7570];
	memory[1892][3] = temp_mem[7571];

	memory[1893][0] = temp_mem[7572];
	memory[1893][1] = temp_mem[7573];
	memory[1893][2] = temp_mem[7574];
	memory[1893][3] = temp_mem[7575];

	memory[1894][0] = temp_mem[7576];
	memory[1894][1] = temp_mem[7577];
	memory[1894][2] = temp_mem[7578];
	memory[1894][3] = temp_mem[7579];

	memory[1895][0] = temp_mem[7580];
	memory[1895][1] = temp_mem[7581];
	memory[1895][2] = temp_mem[7582];
	memory[1895][3] = temp_mem[7583];

	memory[1896][0] = temp_mem[7584];
	memory[1896][1] = temp_mem[7585];
	memory[1896][2] = temp_mem[7586];
	memory[1896][3] = temp_mem[7587];

	memory[1897][0] = temp_mem[7588];
	memory[1897][1] = temp_mem[7589];
	memory[1897][2] = temp_mem[7590];
	memory[1897][3] = temp_mem[7591];

	memory[1898][0] = temp_mem[7592];
	memory[1898][1] = temp_mem[7593];
	memory[1898][2] = temp_mem[7594];
	memory[1898][3] = temp_mem[7595];

	memory[1899][0] = temp_mem[7596];
	memory[1899][1] = temp_mem[7597];
	memory[1899][2] = temp_mem[7598];
	memory[1899][3] = temp_mem[7599];

	memory[1900][0] = temp_mem[7600];
	memory[1900][1] = temp_mem[7601];
	memory[1900][2] = temp_mem[7602];
	memory[1900][3] = temp_mem[7603];

	memory[1901][0] = temp_mem[7604];
	memory[1901][1] = temp_mem[7605];
	memory[1901][2] = temp_mem[7606];
	memory[1901][3] = temp_mem[7607];

	memory[1902][0] = temp_mem[7608];
	memory[1902][1] = temp_mem[7609];
	memory[1902][2] = temp_mem[7610];
	memory[1902][3] = temp_mem[7611];

	memory[1903][0] = temp_mem[7612];
	memory[1903][1] = temp_mem[7613];
	memory[1903][2] = temp_mem[7614];
	memory[1903][3] = temp_mem[7615];

	memory[1904][0] = temp_mem[7616];
	memory[1904][1] = temp_mem[7617];
	memory[1904][2] = temp_mem[7618];
	memory[1904][3] = temp_mem[7619];

	memory[1905][0] = temp_mem[7620];
	memory[1905][1] = temp_mem[7621];
	memory[1905][2] = temp_mem[7622];
	memory[1905][3] = temp_mem[7623];

	memory[1906][0] = temp_mem[7624];
	memory[1906][1] = temp_mem[7625];
	memory[1906][2] = temp_mem[7626];
	memory[1906][3] = temp_mem[7627];

	memory[1907][0] = temp_mem[7628];
	memory[1907][1] = temp_mem[7629];
	memory[1907][2] = temp_mem[7630];
	memory[1907][3] = temp_mem[7631];

	memory[1908][0] = temp_mem[7632];
	memory[1908][1] = temp_mem[7633];
	memory[1908][2] = temp_mem[7634];
	memory[1908][3] = temp_mem[7635];

	memory[1909][0] = temp_mem[7636];
	memory[1909][1] = temp_mem[7637];
	memory[1909][2] = temp_mem[7638];
	memory[1909][3] = temp_mem[7639];

	memory[1910][0] = temp_mem[7640];
	memory[1910][1] = temp_mem[7641];
	memory[1910][2] = temp_mem[7642];
	memory[1910][3] = temp_mem[7643];

	memory[1911][0] = temp_mem[7644];
	memory[1911][1] = temp_mem[7645];
	memory[1911][2] = temp_mem[7646];
	memory[1911][3] = temp_mem[7647];

	memory[1912][0] = temp_mem[7648];
	memory[1912][1] = temp_mem[7649];
	memory[1912][2] = temp_mem[7650];
	memory[1912][3] = temp_mem[7651];

	memory[1913][0] = temp_mem[7652];
	memory[1913][1] = temp_mem[7653];
	memory[1913][2] = temp_mem[7654];
	memory[1913][3] = temp_mem[7655];

	memory[1914][0] = temp_mem[7656];
	memory[1914][1] = temp_mem[7657];
	memory[1914][2] = temp_mem[7658];
	memory[1914][3] = temp_mem[7659];

	memory[1915][0] = temp_mem[7660];
	memory[1915][1] = temp_mem[7661];
	memory[1915][2] = temp_mem[7662];
	memory[1915][3] = temp_mem[7663];

	memory[1916][0] = temp_mem[7664];
	memory[1916][1] = temp_mem[7665];
	memory[1916][2] = temp_mem[7666];
	memory[1916][3] = temp_mem[7667];

	memory[1917][0] = temp_mem[7668];
	memory[1917][1] = temp_mem[7669];
	memory[1917][2] = temp_mem[7670];
	memory[1917][3] = temp_mem[7671];

	memory[1918][0] = temp_mem[7672];
	memory[1918][1] = temp_mem[7673];
	memory[1918][2] = temp_mem[7674];
	memory[1918][3] = temp_mem[7675];

	memory[1919][0] = temp_mem[7676];
	memory[1919][1] = temp_mem[7677];
	memory[1919][2] = temp_mem[7678];
	memory[1919][3] = temp_mem[7679];

	memory[1920][0] = temp_mem[7680];
	memory[1920][1] = temp_mem[7681];
	memory[1920][2] = temp_mem[7682];
	memory[1920][3] = temp_mem[7683];

	memory[1921][0] = temp_mem[7684];
	memory[1921][1] = temp_mem[7685];
	memory[1921][2] = temp_mem[7686];
	memory[1921][3] = temp_mem[7687];

	memory[1922][0] = temp_mem[7688];
	memory[1922][1] = temp_mem[7689];
	memory[1922][2] = temp_mem[7690];
	memory[1922][3] = temp_mem[7691];

	memory[1923][0] = temp_mem[7692];
	memory[1923][1] = temp_mem[7693];
	memory[1923][2] = temp_mem[7694];
	memory[1923][3] = temp_mem[7695];

	memory[1924][0] = temp_mem[7696];
	memory[1924][1] = temp_mem[7697];
	memory[1924][2] = temp_mem[7698];
	memory[1924][3] = temp_mem[7699];

	memory[1925][0] = temp_mem[7700];
	memory[1925][1] = temp_mem[7701];
	memory[1925][2] = temp_mem[7702];
	memory[1925][3] = temp_mem[7703];

	memory[1926][0] = temp_mem[7704];
	memory[1926][1] = temp_mem[7705];
	memory[1926][2] = temp_mem[7706];
	memory[1926][3] = temp_mem[7707];

	memory[1927][0] = temp_mem[7708];
	memory[1927][1] = temp_mem[7709];
	memory[1927][2] = temp_mem[7710];
	memory[1927][3] = temp_mem[7711];

	memory[1928][0] = temp_mem[7712];
	memory[1928][1] = temp_mem[7713];
	memory[1928][2] = temp_mem[7714];
	memory[1928][3] = temp_mem[7715];

	memory[1929][0] = temp_mem[7716];
	memory[1929][1] = temp_mem[7717];
	memory[1929][2] = temp_mem[7718];
	memory[1929][3] = temp_mem[7719];

	memory[1930][0] = temp_mem[7720];
	memory[1930][1] = temp_mem[7721];
	memory[1930][2] = temp_mem[7722];
	memory[1930][3] = temp_mem[7723];

	memory[1931][0] = temp_mem[7724];
	memory[1931][1] = temp_mem[7725];
	memory[1931][2] = temp_mem[7726];
	memory[1931][3] = temp_mem[7727];

	memory[1932][0] = temp_mem[7728];
	memory[1932][1] = temp_mem[7729];
	memory[1932][2] = temp_mem[7730];
	memory[1932][3] = temp_mem[7731];

	memory[1933][0] = temp_mem[7732];
	memory[1933][1] = temp_mem[7733];
	memory[1933][2] = temp_mem[7734];
	memory[1933][3] = temp_mem[7735];

	memory[1934][0] = temp_mem[7736];
	memory[1934][1] = temp_mem[7737];
	memory[1934][2] = temp_mem[7738];
	memory[1934][3] = temp_mem[7739];

	memory[1935][0] = temp_mem[7740];
	memory[1935][1] = temp_mem[7741];
	memory[1935][2] = temp_mem[7742];
	memory[1935][3] = temp_mem[7743];

	memory[1936][0] = temp_mem[7744];
	memory[1936][1] = temp_mem[7745];
	memory[1936][2] = temp_mem[7746];
	memory[1936][3] = temp_mem[7747];

	memory[1937][0] = temp_mem[7748];
	memory[1937][1] = temp_mem[7749];
	memory[1937][2] = temp_mem[7750];
	memory[1937][3] = temp_mem[7751];

	memory[1938][0] = temp_mem[7752];
	memory[1938][1] = temp_mem[7753];
	memory[1938][2] = temp_mem[7754];
	memory[1938][3] = temp_mem[7755];

	memory[1939][0] = temp_mem[7756];
	memory[1939][1] = temp_mem[7757];
	memory[1939][2] = temp_mem[7758];
	memory[1939][3] = temp_mem[7759];

	memory[1940][0] = temp_mem[7760];
	memory[1940][1] = temp_mem[7761];
	memory[1940][2] = temp_mem[7762];
	memory[1940][3] = temp_mem[7763];

	memory[1941][0] = temp_mem[7764];
	memory[1941][1] = temp_mem[7765];
	memory[1941][2] = temp_mem[7766];
	memory[1941][3] = temp_mem[7767];

	memory[1942][0] = temp_mem[7768];
	memory[1942][1] = temp_mem[7769];
	memory[1942][2] = temp_mem[7770];
	memory[1942][3] = temp_mem[7771];

	memory[1943][0] = temp_mem[7772];
	memory[1943][1] = temp_mem[7773];
	memory[1943][2] = temp_mem[7774];
	memory[1943][3] = temp_mem[7775];

	memory[1944][0] = temp_mem[7776];
	memory[1944][1] = temp_mem[7777];
	memory[1944][2] = temp_mem[7778];
	memory[1944][3] = temp_mem[7779];

	memory[1945][0] = temp_mem[7780];
	memory[1945][1] = temp_mem[7781];
	memory[1945][2] = temp_mem[7782];
	memory[1945][3] = temp_mem[7783];

	memory[1946][0] = temp_mem[7784];
	memory[1946][1] = temp_mem[7785];
	memory[1946][2] = temp_mem[7786];
	memory[1946][3] = temp_mem[7787];

	memory[1947][0] = temp_mem[7788];
	memory[1947][1] = temp_mem[7789];
	memory[1947][2] = temp_mem[7790];
	memory[1947][3] = temp_mem[7791];

	memory[1948][0] = temp_mem[7792];
	memory[1948][1] = temp_mem[7793];
	memory[1948][2] = temp_mem[7794];
	memory[1948][3] = temp_mem[7795];

	memory[1949][0] = temp_mem[7796];
	memory[1949][1] = temp_mem[7797];
	memory[1949][2] = temp_mem[7798];
	memory[1949][3] = temp_mem[7799];

	memory[1950][0] = temp_mem[7800];
	memory[1950][1] = temp_mem[7801];
	memory[1950][2] = temp_mem[7802];
	memory[1950][3] = temp_mem[7803];

	memory[1951][0] = temp_mem[7804];
	memory[1951][1] = temp_mem[7805];
	memory[1951][2] = temp_mem[7806];
	memory[1951][3] = temp_mem[7807];

	memory[1952][0] = temp_mem[7808];
	memory[1952][1] = temp_mem[7809];
	memory[1952][2] = temp_mem[7810];
	memory[1952][3] = temp_mem[7811];

	memory[1953][0] = temp_mem[7812];
	memory[1953][1] = temp_mem[7813];
	memory[1953][2] = temp_mem[7814];
	memory[1953][3] = temp_mem[7815];

	memory[1954][0] = temp_mem[7816];
	memory[1954][1] = temp_mem[7817];
	memory[1954][2] = temp_mem[7818];
	memory[1954][3] = temp_mem[7819];

	memory[1955][0] = temp_mem[7820];
	memory[1955][1] = temp_mem[7821];
	memory[1955][2] = temp_mem[7822];
	memory[1955][3] = temp_mem[7823];

	memory[1956][0] = temp_mem[7824];
	memory[1956][1] = temp_mem[7825];
	memory[1956][2] = temp_mem[7826];
	memory[1956][3] = temp_mem[7827];

	memory[1957][0] = temp_mem[7828];
	memory[1957][1] = temp_mem[7829];
	memory[1957][2] = temp_mem[7830];
	memory[1957][3] = temp_mem[7831];

	memory[1958][0] = temp_mem[7832];
	memory[1958][1] = temp_mem[7833];
	memory[1958][2] = temp_mem[7834];
	memory[1958][3] = temp_mem[7835];

	memory[1959][0] = temp_mem[7836];
	memory[1959][1] = temp_mem[7837];
	memory[1959][2] = temp_mem[7838];
	memory[1959][3] = temp_mem[7839];

	memory[1960][0] = temp_mem[7840];
	memory[1960][1] = temp_mem[7841];
	memory[1960][2] = temp_mem[7842];
	memory[1960][3] = temp_mem[7843];

	memory[1961][0] = temp_mem[7844];
	memory[1961][1] = temp_mem[7845];
	memory[1961][2] = temp_mem[7846];
	memory[1961][3] = temp_mem[7847];

	memory[1962][0] = temp_mem[7848];
	memory[1962][1] = temp_mem[7849];
	memory[1962][2] = temp_mem[7850];
	memory[1962][3] = temp_mem[7851];

	memory[1963][0] = temp_mem[7852];
	memory[1963][1] = temp_mem[7853];
	memory[1963][2] = temp_mem[7854];
	memory[1963][3] = temp_mem[7855];

	memory[1964][0] = temp_mem[7856];
	memory[1964][1] = temp_mem[7857];
	memory[1964][2] = temp_mem[7858];
	memory[1964][3] = temp_mem[7859];

	memory[1965][0] = temp_mem[7860];
	memory[1965][1] = temp_mem[7861];
	memory[1965][2] = temp_mem[7862];
	memory[1965][3] = temp_mem[7863];

	memory[1966][0] = temp_mem[7864];
	memory[1966][1] = temp_mem[7865];
	memory[1966][2] = temp_mem[7866];
	memory[1966][3] = temp_mem[7867];

	memory[1967][0] = temp_mem[7868];
	memory[1967][1] = temp_mem[7869];
	memory[1967][2] = temp_mem[7870];
	memory[1967][3] = temp_mem[7871];

	memory[1968][0] = temp_mem[7872];
	memory[1968][1] = temp_mem[7873];
	memory[1968][2] = temp_mem[7874];
	memory[1968][3] = temp_mem[7875];

	memory[1969][0] = temp_mem[7876];
	memory[1969][1] = temp_mem[7877];
	memory[1969][2] = temp_mem[7878];
	memory[1969][3] = temp_mem[7879];

	memory[1970][0] = temp_mem[7880];
	memory[1970][1] = temp_mem[7881];
	memory[1970][2] = temp_mem[7882];
	memory[1970][3] = temp_mem[7883];

	memory[1971][0] = temp_mem[7884];
	memory[1971][1] = temp_mem[7885];
	memory[1971][2] = temp_mem[7886];
	memory[1971][3] = temp_mem[7887];

	memory[1972][0] = temp_mem[7888];
	memory[1972][1] = temp_mem[7889];
	memory[1972][2] = temp_mem[7890];
	memory[1972][3] = temp_mem[7891];

	memory[1973][0] = temp_mem[7892];
	memory[1973][1] = temp_mem[7893];
	memory[1973][2] = temp_mem[7894];
	memory[1973][3] = temp_mem[7895];

	memory[1974][0] = temp_mem[7896];
	memory[1974][1] = temp_mem[7897];
	memory[1974][2] = temp_mem[7898];
	memory[1974][3] = temp_mem[7899];

	memory[1975][0] = temp_mem[7900];
	memory[1975][1] = temp_mem[7901];
	memory[1975][2] = temp_mem[7902];
	memory[1975][3] = temp_mem[7903];

	memory[1976][0] = temp_mem[7904];
	memory[1976][1] = temp_mem[7905];
	memory[1976][2] = temp_mem[7906];
	memory[1976][3] = temp_mem[7907];

	memory[1977][0] = temp_mem[7908];
	memory[1977][1] = temp_mem[7909];
	memory[1977][2] = temp_mem[7910];
	memory[1977][3] = temp_mem[7911];

	memory[1978][0] = temp_mem[7912];
	memory[1978][1] = temp_mem[7913];
	memory[1978][2] = temp_mem[7914];
	memory[1978][3] = temp_mem[7915];

	memory[1979][0] = temp_mem[7916];
	memory[1979][1] = temp_mem[7917];
	memory[1979][2] = temp_mem[7918];
	memory[1979][3] = temp_mem[7919];

	memory[1980][0] = temp_mem[7920];
	memory[1980][1] = temp_mem[7921];
	memory[1980][2] = temp_mem[7922];
	memory[1980][3] = temp_mem[7923];

	memory[1981][0] = temp_mem[7924];
	memory[1981][1] = temp_mem[7925];
	memory[1981][2] = temp_mem[7926];
	memory[1981][3] = temp_mem[7927];

	memory[1982][0] = temp_mem[7928];
	memory[1982][1] = temp_mem[7929];
	memory[1982][2] = temp_mem[7930];
	memory[1982][3] = temp_mem[7931];

	memory[1983][0] = temp_mem[7932];
	memory[1983][1] = temp_mem[7933];
	memory[1983][2] = temp_mem[7934];
	memory[1983][3] = temp_mem[7935];

	memory[1984][0] = temp_mem[7936];
	memory[1984][1] = temp_mem[7937];
	memory[1984][2] = temp_mem[7938];
	memory[1984][3] = temp_mem[7939];

	memory[1985][0] = temp_mem[7940];
	memory[1985][1] = temp_mem[7941];
	memory[1985][2] = temp_mem[7942];
	memory[1985][3] = temp_mem[7943];

	memory[1986][0] = temp_mem[7944];
	memory[1986][1] = temp_mem[7945];
	memory[1986][2] = temp_mem[7946];
	memory[1986][3] = temp_mem[7947];

	memory[1987][0] = temp_mem[7948];
	memory[1987][1] = temp_mem[7949];
	memory[1987][2] = temp_mem[7950];
	memory[1987][3] = temp_mem[7951];

	memory[1988][0] = temp_mem[7952];
	memory[1988][1] = temp_mem[7953];
	memory[1988][2] = temp_mem[7954];
	memory[1988][3] = temp_mem[7955];

	memory[1989][0] = temp_mem[7956];
	memory[1989][1] = temp_mem[7957];
	memory[1989][2] = temp_mem[7958];
	memory[1989][3] = temp_mem[7959];

	memory[1990][0] = temp_mem[7960];
	memory[1990][1] = temp_mem[7961];
	memory[1990][2] = temp_mem[7962];
	memory[1990][3] = temp_mem[7963];

	memory[1991][0] = temp_mem[7964];
	memory[1991][1] = temp_mem[7965];
	memory[1991][2] = temp_mem[7966];
	memory[1991][3] = temp_mem[7967];

	memory[1992][0] = temp_mem[7968];
	memory[1992][1] = temp_mem[7969];
	memory[1992][2] = temp_mem[7970];
	memory[1992][3] = temp_mem[7971];

	memory[1993][0] = temp_mem[7972];
	memory[1993][1] = temp_mem[7973];
	memory[1993][2] = temp_mem[7974];
	memory[1993][3] = temp_mem[7975];

	memory[1994][0] = temp_mem[7976];
	memory[1994][1] = temp_mem[7977];
	memory[1994][2] = temp_mem[7978];
	memory[1994][3] = temp_mem[7979];

	memory[1995][0] = temp_mem[7980];
	memory[1995][1] = temp_mem[7981];
	memory[1995][2] = temp_mem[7982];
	memory[1995][3] = temp_mem[7983];

	memory[1996][0] = temp_mem[7984];
	memory[1996][1] = temp_mem[7985];
	memory[1996][2] = temp_mem[7986];
	memory[1996][3] = temp_mem[7987];

	memory[1997][0] = temp_mem[7988];
	memory[1997][1] = temp_mem[7989];
	memory[1997][2] = temp_mem[7990];
	memory[1997][3] = temp_mem[7991];

	memory[1998][0] = temp_mem[7992];
	memory[1998][1] = temp_mem[7993];
	memory[1998][2] = temp_mem[7994];
	memory[1998][3] = temp_mem[7995];

	memory[1999][0] = temp_mem[7996];
	memory[1999][1] = temp_mem[7997];
	memory[1999][2] = temp_mem[7998];
	memory[1999][3] = temp_mem[7999];

end

assign o_instr = memory[i_pc[31:2]];

endmodule
